*  
* Diode Model Produced by Altium Ltd  
* Date:  10-Mar-2004 
*  
* Manufacturer: Agilent  
* Component Name: HDSP-F153  
*  
* Parameters derived from information available in data sheet.  
*  
*                 common-cathode 
*                 |  anode-f 
*                 |  |  anode-g 
*                 |  |  |  anode-e 
*                 |  |  |  |  anode-d 
*                 |  |  |  |  |  common-cathode 
*                 |  |  |  |  |  |  anode-DP 
*                 |  |  |  |  |  |  |  anode-c 
*                 |  |  |  |  |  |  |  |  anode-b 
*                 |  |  |  |  |  |  |  |  |  anode-a
*                 |  |  |  |  |  |  |  |  |  |
.SUBCKT HDSP_F153 1  2  3  4  5  6  7  8  9  10

DA1  10 1 dHDSP_F153
DB1   9 1 dHDSP_F153
DC1   8 1 dHDSP_F153
DD1   5 1 dHDSP_F153
DE1   4 1 dHDSP_F153
DF1   2 1 dHDSP_F153
DG1   3 1 dHDSP_F153
DDP1  7 1 dHDSP_F153

DA2  10 6 dHDSP_F153
DB2   9 6 dHDSP_F153
DC2   8 6 dHDSP_F153
DD2   5 6 dHDSP_F153
DE2   4 6 dHDSP_F153
DF2   2 6 dHDSP_F153
DG2   3 6 dHDSP_F153
DDP2  7 6 dHDSP_F153

.MODEL dHDSP_F153 D
+ (  
+    IS  = 1.31055154E-15 
+     N  = 2.20660855 
+    RS  = 1.60736539 
+    BV  = 14.25
+   IBV  = 100u
+ )  

.ENDS HDSP_F153
*  
* Diode Model Produced by Altium Ltd  
* Date:  10-Mar-2004 
*  
* Manufacturer: Agilent  
* Component Name: HDSP-303A  
*  
* Parameters derived from information available in data sheet.  
*
*                 anode-G
*                 |  anode-F
*                 |  |  comon-cathode
*                 |  |  |  anode-E
*                 |  |  |  |  anode-D
*                 |  |  |  |  |  anode-DP
*                 |  |  |  |  |  |  anode-C
*                 |  |  |  |  |  |  |  comon-cathode
*                 |  |  |  |  |  |  |  |  anode-B
*                 |  |  |  |  |  |  |  |  |  anode-A
*                 |  |  |  |  |  |  |  |  |  |  
.SUBCKT HDSP_303A 1  2  3  4  5  6  7  8  9  10

DA1  10  3  dHDSP_303A
DB1   9  3  dHDSP_303A
DC1   7  3  dHDSP_303A
DD1   5  3  dHDSP_303A
DE1   4  3  dHDSP_303A
DF1   2  3  dHDSP_303A
DG1   1  3  dHDSP_303A
DDP1  6  3  dHDSP_303A

DA2  10  8  dHDSP_303A
DB2   9  8  dHDSP_303A
DC2   7  8  dHDSP_303A
DD2   5  8  dHDSP_303A
DE2   4  8  dHDSP_303A
DF2   2  8  dHDSP_303A
DG2   1  8  dHDSP_303A
DDP2  6  8  dHDSP_303A

.MODEL dHDSP_303A D
+ (  
+    IS = 4.59961571E-15 
+     N = 2.40621673 
+    RS = 1.90931135 
+    BV = 4.5
+   IBV = 100u
+ )  

.ENDS HDSP_303A
*  
* Diode Model Produced by Altium Ltd  
* Date:  10-Mar-2004 
*  
* Manufacturer: Agilent  
* Component Name: HDSP-563G  
*  
* Parameters derived from information available in data sheet.  
*
*                 anode-E
*                 |  anode-D
*                 |  |  comon-cathode
*                 |  |  |  anode-C
*                 |  |  |  |  anode-DP
*                 |  |  |  |  |  anode-B
*                 |  |  |  |  |  |  anode-A
*                 |  |  |  |  |  |  |  comon-cathode
*                 |  |  |  |  |  |  |  |  anode-F
*                 |  |  |  |  |  |  |  |  |  anode-G
*                 |  |  |  |  |  |  |  |  |  |  
.SUBCKT HDSP_563G 1  2  3  4  5  6  7  8  9  10

DA1   7  3  dHDSP_563G
DB1   6  3  dHDSP_563G
DC1   4  3  dHDSP_563G
DD1   2  3  dHDSP_563G
DE1   1  3  dHDSP_563G
DF1   9  3  dHDSP_563G
DG1  10  3  dHDSP_563G
DDP1  5  3  dHDSP_563G

DA2   7  8  dHDSP_563G
DB2   6  8  dHDSP_563G
DC2   4  8  dHDSP_563G
DD2   2  8  dHDSP_563G
DE2   1  8  dHDSP_563G
DF2   9  8  dHDSP_563G
DG2  10  8  dHDSP_563G
DDP2  5  8  dHDSP_563G

.MODEL dHDSP_563G D
+ (  
+     IS = 3.14401041E-29 
+      N = 1.25233679 
+     RS = 9.99993505 
+     BV = 4.8 
+    IBV = 100u 
+ )  

.ENDS HDSP_563G
*  
* Diode Model Produced by Altium Ltd  
* Date:  10-Mar-2004 
*  
* Manufacturer: Agilent  
* Component Name: HDSP-H513  
*  
* Parameters derived from information available in data sheet.  
* 
*                 anode-e
*                 |  anode-d
*                 |  |  common-cathode
*                 |  |  |  anode-c
*                 |  |  |  |  anode-DP
*                 |  |  |  |  |  anode-b
*                 |  |  |  |  |  |  anode-a
*                 |  |  |  |  |  |  |  common-cathode
*                 |  |  |  |  |  |  |  |  anode-f
*                 |  |  |  |  |  |  |  |  |  anode-g
*                 |  |  |  |  |  |  |  |  |  | 
.SUBCKT HDSP_H513 1  2  3  4  5  6  7  8  9  10

DA1    7  3  dHDSP_H513
DB1    6  3  dHDSP_H513
DC1    4  3  dHDSP_H513
DD1    2  3  dHDSP_H513
DE1    1  3  dHDSP_H513
DF1    9  3  dHDSP_H513
DG1   10  3  dHDSP_H513
DDP1   5  3  dHDSP_H513

DA2    7  8  dHDSP_H513
DB2    6  8  dHDSP_H513
DC2    4  8  dHDSP_H513
DD2    2  8  dHDSP_H513
DE2    1  8  dHDSP_H513
DF2    9  8  dHDSP_H513
DG2   10  8  dHDSP_H513
DDP2   5  8  dHDSP_H513

.MODEL dHDSP_H513 D
+ (  
+     IS = 1.61114016E-27 
+      N = 1.30291189 
+     RS = 12.83456794 
+     BV = 50 
+    IBV = 100u 
+ )  

.ENDS HDSP_H513
*  
* Diode Model Produced by Altium Ltd  
* Date:  10-Mar-2004 
*  
* Manufacturer: Agilent  
* Component Name: HDSP-313G  
*  
* Parameters derived from information available in data sheet.  
*  
*                 anode-G 
*                 |  anode-F 
*                 |  |  common-cathode 
*                 |  |  |  anode-E 
*                 |  |  |  |  anode-D 
*                 |  |  |  |  |  anode-DP 
*                 |  |  |  |  |  |  anode-C 
*                 |  |  |  |  |  |  |  common-cathode 
*                 |  |  |  |  |  |  |  |  anode-B 
*                 |  |  |  |  |  |  |  |  |  anode-A
*                 |  |  |  |  |  |  |  |  |  |
.SUBCKT HDSP_313G 1  2  3  4  5  6  7  8  9  10

DA1  3  10 dHDSP_313G
DB1  3   9 dHDSP_313G
DC1  3   7 dHDSP_313G
DD1  3   5 dHDSP_313G
DE1  3   4 dHDSP_313G
DF1  3   2 dHDSP_313G
DG1  3   1 dHDSP_313G
DDP1 3   6 dHDSP_313G

DA2  8  10 dHDSP_313G
DB2  8   9 dHDSP_313G
DC2  8   7 dHDSP_313G
DD2  8   5 dHDSP_313G
DE2  8   4 dHDSP_313G
DF2  8   2 dHDSP_313G
DG2  8   1 dHDSP_313G
DDP2 8   6 dHDSP_313G

.MODEL dHDSP_313G D
+ (  
+     IS = 1.61114016E-27 
+      N = 1.30291189 
+     RS = 12.83456794 
+     BV = 50 
+    IBV = 100u 
+ )  

.ENDS HDSP_313G
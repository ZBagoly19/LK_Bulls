*  
* Diode Model Produced by Altium Ltd  
* Date:  3-May-2004 
*  
* Manufacturer: Renesas  
* Component Name: HDSP-A403  
*  
* Parameters derived from information available in data sheet.  
* 
*                 common-cathode
*                 |  anode-f
*                 |  |  anode-g
*                 |  |  |  anode-e
*                 |  |  |  |  anode-d
*                 |  |  |  |  |  common-cathode
*                 |  |  |  |  |  |  anode-DP
*                 |  |  |  |  |  |  |  anode-c
*                 |  |  |  |  |  |  |  |  anode-b
*                 |  |  |  |  |  |  |  |  |  anode-a
*                 |  |  |  |  |  |  |  |  |  |
.SUBCKT HDSP_A403 1  2  3  4  5  6  7  8  9  10

DA1  10  1  dHDSP_A403
DB1   9  1  dHDSP_A403
DC1   8  1  dHDSP_A403
DD1   5  1  dHDSP_A403
DE1   4  1  dHDSP_A403
DF1   2  1  dHDSP_A403
DG1   3  1  dHDSP_A403
DDP1  7  1  dHDSP_A403

DA2  10  6  dHDSP_A403
DB2   9  6  dHDSP_A403
DC2   8  6  dHDSP_A403
DD2   5  6  dHDSP_A403
DE2   4  6  dHDSP_A403
DF2   2  6  dHDSP_A403
DG2   3  6  dHDSP_A403
DDP2  7  6  dHDSP_A403

.MODEL dHDSP_A403 D
+ (  
+     IS = 1.31238168E-27 
+      N = 1.06196807 
+     RS = 24.48189481 
+     BV = 25
+    IBV = 100u 
+ ) 

.ENDS HDSP_A403
*  
* Diode Model Produced by Altium Ltd  
* Date:  3-May-2004 
*  
* Manufacturer: Renesas  
* Component Name: HDSP-7501  
*  
* Parameters derived from information available in data sheet.  
* 
*                 common-anode
*                 |  cathode-f
*                 |  |  cathode-g
*                 |  |  |  cathode-e
*                 |  |  |  |  cathode-d
*                 |  |  |  |  |  common-anode
*                 |  |  |  |  |  |  cathode-DP
*                 |  |  |  |  |  |  |  cathode-c
*                 |  |  |  |  |  |  |  |  cathode-b
*                 |  |  |  |  |  |  |  |  |  cathode-a
*                 |  |  |  |  |  |  |  |  |  |
.SUBCKT HDSP_7501 1  2  3  4  5  6  7  8  9  10

DA1  1  10  dHDSP_7501
DB1  1   9  dHDSP_7501
DC1  1   8  dHDSP_7501
DD1  1   5  dHDSP_7501
DE1  1   4  dHDSP_7501
DF1  1   2  dHDSP_7501
DG1  1   3  dHDSP_7501
DDP1 1   7  dHDSP_7501

DA2  6  10  dHDSP_7501
DB2  6   9  dHDSP_7501
DC2  6   8  dHDSP_7501
DD2  6   5  dHDSP_7501
DE2  6   4  dHDSP_7501
DF2  6   2  dHDSP_7501
DG2  6   3  dHDSP_7501
DDP2 6   7  dHDSP_7501

.MODEL dHDSP_7501 D
+ (  
+     IS = 1.31238168E-27 
+      N = 1.06196807 
+     RS = 24.48189481 
+     BV = 25
+    IBV = 100u 
+ )  

.ENDS HDSP_7501
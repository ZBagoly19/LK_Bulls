*  
* Diode Model Produced by Altium Ltd  
* Date:  10-Mar-2004 
*  
* Manufacturer: Agilent  
* Component Name: HDSP-U503  
*  
* Parameters derived from information available in data sheet.  
*  
*                  anode-a 
*                  |  anode-f 
*                  |  |  anode-g 
*                  |  |  |  anode-e 
*                  |  |  |  |  anode-d 
*                  |  |  |  |  |  cathode-DP 
*                  |  |  |  |  |  |  anode-DP 
*                  |  |  |  |  |  |  |  anode-c 
*                  |  |  |  |  |  |  |  |  common-cathode 
*                  |  |  |  |  |  |  |  |  |  anode-b
*                  |  |  |  |  |  |  |  |  |  |
.SUBCKT HDSP_U503 1  2  3  4  5  6  7  8  9  10

D1  1  9 dHDSP_U503
D2  2  9 dHDSP_U503
D3  3  9 dHDSP_U503
D4  4  9 dHDSP_U503
D5  5  9 dHDSP_U503
D6  7  6 dHDSP_U503
D7  8  9 dHDSP_U503
D8 10  9 dHDSP_U503

.MODEL dHDSP_U503 D
+ (  
+     IS = 1.61114016E-27 
+      N = 1.30291189 
+     RS = 12.83456794 
+     BV = 50 
+    IBV = 100u 
+ )  

.ENDS HDSP_U503
*  
* Diode Model Produced by Altium Ltd  
* Date:  11-Mar-2004 
*  
* Manufacturer: Agilent  
* Component Name: HDSP-563C  
*  
* Parameters derived from information available in data sheet.  
* 
*                 anode-e
*                 |  anode-d
*                 |  |  common-cathode
*                 |  |  |  anode-c
*                 |  |  |  |  anode-DP
*                 |  |  |  |  |  anode-b
*                 |  |  |  |  |  |  anode-a
*                 |  |  |  |  |  |  |  common-cathode
*                 |  |  |  |  |  |  |  |  anode-f
*                 |  |  |  |  |  |  |  |  |  anode-g
*                 |  |  |  |  |  |  |  |  |  |
.SUBCKT HDSP_563C 1  2  3  4  5  6  7  8  9  10

DA1   7  3 dHDSP_563C
DB1   6  3 dHDSP_563C
DC1   4  3 dHDSP_563C
DD1   2  3 dHDSP_563C
DE1   1  3 dHDSP_563C
DF1   9  3 dHDSP_563C
DG1  10  3 dHDSP_563C
DDP1  5  3 dHDSP_563C

DA2   7  8 dHDSP_563C
DB2   6  8 dHDSP_563C
DC2   4  8 dHDSP_563C
DD2   2  8 dHDSP_563C
DE2   1  8 dHDSP_563C
DF2   9  8 dHDSP_563C
DG2  10  8 dHDSP_563C
DDP2  5  8 dHDSP_563C

 
.MODEL dHDSP_563C D
+ (  
+    IS = 2.34165185E-18 
+     N = 1.64080796 
+    RS = 5.35791037 
+    BV = 4.5
+   IBV = 100u
+ )  

.ENDS HDSP_563C
*  
* Diode Model Produced by Altium Ltd  
* Date:  7-Apr-2004 
*  
* Manufacturer: Agilent  
* Component Name: HDSP-515H  
*  
* Parameters derived from information available in data sheet.  
* 
*                 e - cathode
*                 |  d - cathode
*                 |  |  common-anode
*                 |  |  |  c - cathode
*                 |  |  |  |  DP - cathode
*                 |  |  |  |  |  b - cathode
*                 |  |  |  |  |  |  a - cathode
*                 |  |  |  |  |  |  |  common-anode
*                 |  |  |  |  |  |  |  |  f - cathode
*                 |  |  |  |  |  |  |  |  |  g - cathode
*                 |  |  |  |  |  |  |  |  |  | 
.SUBCKT HDSP_515H 1  2  3  4  5  6  7  8  9  10

DA1  3  7 dHDSP_515H
DB1  3  6 dHDSP_515H
DC1  3  4 dHDSP_515H
DD1  3  2 dHDSP_515H
DE1  3  1 dHDSP_515H
DF1  3  9 dHDSP_515H
DG1  3 10 dHDSP_515H
DDP1 3  5 dHDSP_515H

DA2  8  7 dHDSP_515H
DB2  8  6 dHDSP_515H
DC2  8  4 dHDSP_515H
DD2  8  2 dHDSP_515H
DE2  8  1 dHDSP_515H
DF2  8  9 dHDSP_515H
DG2  8 10 dHDSP_515H
DDP2 8  5 dHDSP_515H

.MODEL dHDSP_515H D
+ (  
+    IS  = 2.08276754E-16 
+     N  = 2.17799178 
+    RS  = 0.50892350
+    BV  = 14.25
+   IBV  = 100u
+ )  

.ENDS HDSP_515H
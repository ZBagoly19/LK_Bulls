*  
* Diode Model Produced by Altium Ltd  
* Date:  10-Mar-2004 
*  
* Manufacturer: Agilent  
* Component Name: HDSP-561A  
*  
* Parameters derived from information available in data sheet.  
*
*                 cathode-E
*                 |  cathode-D
*                 |  |  comon-anode
*                 |  |  |  cathode-C
*                 |  |  |  |  cathode-DP
*                 |  |  |  |  |  cathode-B
*                 |  |  |  |  |  |  cathode-A
*                 |  |  |  |  |  |  |  comon-anode
*                 |  |  |  |  |  |  |  |  cathode-F
*                 |  |  |  |  |  |  |  |  |  cathode-G
*                 |  |  |  |  |  |  |  |  |  |  
.SUBCKT HDSP_561A 1  2  3  4  5  6  7  8  9  10

DA1  3   7 dHDSP_561A
DB1  3   6 dHDSP_561A
DC1  3   4 dHDSP_561A
DD1  3   2 dHDSP_561A
DE1  3   1 dHDSP_561A
DF1  3   9 dHDSP_561A
DG1  3  10 dHDSP_561A
DDP1 3   5 dHDSP_561A

DA2  8   7 dHDSP_561A
DB2  8   6 dHDSP_561A
DC2  8   4 dHDSP_561A
DD2  8   2 dHDSP_561A
DE2  8   1 dHDSP_561A
DF2  8   9 dHDSP_561A
DG2  8  10 dHDSP_561A
DDP2 8   5 dHDSP_561A

.MODEL dHDSP_561A D
+ (  
+    IS = 4.59961571E-15 
+     N = 2.40621673 
+    RS = 1.90931135 
+    BV = 4.5
+   IBV = 100u
+ )  

.ENDS HDSP_561A
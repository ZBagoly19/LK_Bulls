*  
* Diode Model Produced by Altium Ltd  
* Date:  7-Apr-2004 
*  
* Manufacturer: Agilent  
* Component Name: HDSP-H103  
*  
* Parameters derived from information available in data sheet.  
* 
*                 anode-e
*                 |  anode-d
*                 |  |  common-cathode
*                 |  |  |  anode-c
*                 |  |  |  |  anode-DP
*                 |  |  |  |  |  anode-b
*                 |  |  |  |  |  |  anode-a
*                 |  |  |  |  |  |  |  common-cathode
*                 |  |  |  |  |  |  |  |  anode-f
*                 |  |  |  |  |  |  |  |  |  anode-g
*                 |  |  |  |  |  |  |  |  |  |  
.SUBCKT HDSP_H103 1  2  3  4  5  6  7  8  9  10

DA1   7  3  dHDSP_H103
DB1   6  3  dHDSP_H103
DC1   4  3  dHDSP_H103
DD1   2  3  dHDSP_H103
DE1   1  3  dHDSP_H103
DF1   9  3  dHDSP_H103
DG1  10  3  dHDSP_H103
DDP1  5  3  dHDSP_H103

DA2   7  8  dHDSP_H103
DB2   6  8  dHDSP_H103
DC2   4  8  dHDSP_H103
DD2   2  8  dHDSP_H103
DE2   1  8  dHDSP_H103
DF2   9  8  dHDSP_H103
DG2  10  8  dHDSP_H103
DDP2  5  8  dHDSP_H103

.MODEL dHDSP_H103 D
+ (  
+    IS  = 2.08276754E-16 
+     N  = 2.17799178 
+    RS  = 0.50892350
+    BV  = 14.25
+   IBV  = 100u
+ )  

.ENDS HDSP_H103
*  
* Diode Model Produced by Altium Ltd  
* Date:  10-Mar-2004 
*  
* Manufacturer: Agilent  
* Component Name: HDSP-301A  
*  
* Parameters derived from information available in data sheet.  
*
*                 cathode-G
*                 |  cathode-F
*                 |  |  comon-anode
*                 |  |  |  cathode-E
*                 |  |  |  |  cathode-D
*                 |  |  |  |  |  cathode-DP
*                 |  |  |  |  |  |  cathode-C
*                 |  |  |  |  |  |  |  comon-anode
*                 |  |  |  |  |  |  |  |  cathode-B
*                 |  |  |  |  |  |  |  |  |  cathode-A
*                 |  |  |  |  |  |  |  |  |  |  
.SUBCKT HDSP_301A 1  2  3  4  5  6  7  8  9  10

DA1  3  10 dHDSP_301A
DB1  3   9 dHDSP_301A
DC1  3   7 dHDSP_301A
DD1  3   5 dHDSP_301A
DE1  3   4 dHDSP_301A
DF1  3   2 dHDSP_301A
DG1  3   1 dHDSP_301A
DDP1 3   6 dHDSP_301A

DA2  8  10 dHDSP_301A
DB2  8   9 dHDSP_301A
DC2  8   7 dHDSP_301A
DD2  8   5 dHDSP_301A
DE2  8   4 dHDSP_301A
DF2  8   2 dHDSP_301A
DG2  8   1 dHDSP_301A
DDP2 8   6 dHDSP_301A

.MODEL dHDSP_301A D
+ (  
+    IS = 4.59961571E-15 
+     N = 2.40621673 
+    RS = 1.90931135 
+    BV = 4.5
+   IBV = 100u
+ )  

.ENDS HDSP_301A
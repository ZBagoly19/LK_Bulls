*  
* Diode Model Produced by Altium Ltd  
* Date:  10-Mar-2004 
*  
* Manufacturer: Agilent  
* Component Name: HDSP-N101  
*  
* Parameters derived from information available in data sheet.  
*
*                 cathode-a
*                 |  cathode-f
*                 |  |  common-anode
*                 |  |  |  cathode-e
*                 |  |  |  |  common-anode
*                 |  |  |  |  |  cathode-DP
*                 |  |  |  |  |  |  cathode-d
*                 |  |  |  |  |  |  |  common-anode
*                 |  |  |  |  |  |  |  |  cathode-c
*                 |  |  |  |  |  |  |  |  |  cathode-g
*                 |  |  |  |  |  |  |  |  |  |  cathode-b
*                 |  |  |  |  |  |  |  |  |  |  |  common-anode
*                 |  |  |  |  |  |  |  |  |  |  |  |
.SUBCKT HDSP_N101 2  3  4  5  6  10 11 12 13 14 15 17

DA1   4   2  dHDSP_N101
DB1   4  15  dHDSP_N101
DC1   4  13  dHDSP_N101
DD1   4  11  dHDSP_N101
DE1   4   5  dHDSP_N101
DF1   4   3  dHDSP_N101
DG1   4  14  dHDSP_N101
DDP1  4  10  dHDSP_N101

DA2   6   2  dHDSP_N101
DB2   6  15  dHDSP_N101
DC2   6  13  dHDSP_N101
DD2   6  11  dHDSP_N101
DE2   6   5  dHDSP_N101
DF2   6   3  dHDSP_N101
DG2   6  14  dHDSP_N101
DDP2  6  10  dHDSP_N101

DA3  12    2  dHDSP_N101
DB3  12   15  dHDSP_N101
DC3  12   13  dHDSP_N101
DD3  12   11  dHDSP_N101
DE3  12    5  dHDSP_N101
DF3  12    3  dHDSP_N101
DG3  12   14  dHDSP_N101
DDP3 12   10  dHDSP_N101

DA4  17    2  dHDSP_N101
DB4  17   15  dHDSP_N101
DC4  17   13  dHDSP_N101
DD4  17   11  dHDSP_N101
DE4  17    5  dHDSP_N101
DF4  17    3  dHDSP_N101
DG4  17   14  dHDSP_N101
DDP4 17   10  dHDSP_N101
  
.MODEL dHDSP_N101 D
+ (  
+    IS  = 2.08276754E-16 
+     N  = 2.17799178 
+    RS  = 0.50892350
+    BV  = 14.25
+   IBV  = 100u
+ )  

.ENDS HDSP_N101
*  
* Diode Model Produced by Altium Ltd  
* Date:  7-Apr-2004 
*  
* Manufacturer: Agilent  
* Component Name: HDSP-816E  
*  
* Parameters derived from information available in data sheet.  
*  
*                 anode-a
*                 |  anode-f
*                 |  |  common-cathode
*                 |  |  |  anode-e
*                 |  |  |  |  common-cathode
*                 |  |  |  |  |  anode-DP
*                 |  |  |  |  |  |  anode-d
*                 |  |  |  |  |  |  |  common-cathode
*                 |  |  |  |  |  |  |  |  anode-c
*                 |  |  |  |  |  |  |  |  |  anode-g
*                 |  |  |  |  |  |  |  |  |  |  anode-b
*                 |  |  |  |  |  |  |  |  |  |  |  common-cathode
*                 |  |  |  |  |  |  |  |  |  |  |  |
.SUBCKT HDSP_816E 1  2  3  4  5  9  10 11 12 13 14 16

DA1    1  3  dHDSP_816E
DB1   14  3  dHDSP_816E
DC1   12  3  dHDSP_816E
DD1   10  3  dHDSP_816E
DE1    4  3  dHDSP_816E
DF1    2  3  dHDSP_816E
DG1   13  3  dHDSP_816E
DDP1   9  3  dHDSP_816E

DA2    1  5  dHDSP_816E
DB2   14  5  dHDSP_816E
DC2   12  5  dHDSP_816E
DD2   10  5  dHDSP_816E
DE2    4  5  dHDSP_816E
DF2    2  5  dHDSP_816E
DG2   13  5  dHDSP_816E
DDP2   9  5  dHDSP_816E

DA3    1 11  dHDSP_816E
DB3   14 11  dHDSP_816E
DC3   12 11  dHDSP_816E
DD3   10 11  dHDSP_816E
DE3    4 11  dHDSP_816E
DF3    2 11  dHDSP_816E
DG3   13 11  dHDSP_816E
DDP3   9 11  dHDSP_816E

DA4    1 16  dHDSP_816E
DB4   14 16  dHDSP_816E
DC4   12 16  dHDSP_816E
DD4   10 16  dHDSP_816E
DE4    4 16  dHDSP_816E
DF4    2 16  dHDSP_816E
DG4   13 16  dHDSP_816E
DDP4   9 16  dHDSP_816E

.MODEL dHDSP_816E D
+ (  
+     IS = 1.16713374E-20 
+      N = 1.46891103 
+     RS = 23.91420160 
+     BV = 25
+    IBV = 100u 
+ )  

.ENDS HDSP_816E
*  
* Diode Model Produced by Altium Ltd  
* Date:  7-Apr-2004 
*  
* Manufacturer: Agilent  
* Component Name: 5082-7653  
*  
* Parameters derived from information available in data sheet.  
* 
*                 anode-a
*                 |  anode-f
*                 |  |  common-cathode
*                 |  |  |  anode-e
*                 |  |  |  |  anode-d
*                 |  |  |  |  |  anode-DP
*                 |  |  |  |  |  |  anode-c
*                 |  |  |  |  |  |  |  anode-g
*                 |  |  |  |  |  |  |  |  anode-b
*                 |  |  |  |  |  |  |  |  |  common-cathode
*                 |  |  |  |  |  |  |  |  |  |
.SUBCKT 5082_7653 1  2  3  7  8  9  10 11 13 14

DA1   1  3 d5082_7653
DB1  13  3 d5082_7653
DC1  10  3 d5082_7653
DD1   8  3 d5082_7653
DE1   7  3 d5082_7653
DF1   2  3 d5082_7653
DG1  11  3 d5082_7653
DDP1  9  3 d5082_7653

DA2   1 14 d5082_7653
DB2  13 14 d5082_7653
DC2  10 14 d5082_7653
DD2   8 14 d5082_7653
DE2   7 14 d5082_7653
DF2   2 14 d5082_7653
DG2  11 14 d5082_7653
DDP2  9 14 d5082_7653

.MODEL d5082_7653 D
+ (  
+     IS = 1.95991353E-12 
+      N = 2.90687588 
+     RS = 18.38470387 
+     BV = 30
+    IBV = 100u 
+ )  

.ENDS 5082_7653
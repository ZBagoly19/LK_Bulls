*  
* Diode Model Produced by Altium Ltd  
* Date:  6-Apr-2004 
*  
* Manufacturer: Agilent  
* Component Name: HDSP-H403  
*  
* Parameters derived from information available in data sheet.  
* 
*                 anode-e
*                 |  anode-d
*                 |  |  common-cathode
*                 |  |  |  anode-c
*                 |  |  |  |  anode-DP
*                 |  |  |  |  |  anode-b
*                 |  |  |  |  |  |  anode-a
*                 |  |  |  |  |  |  |  common-cathode
*                 |  |  |  |  |  |  |  |  anode-f
*                 |  |  |  |  |  |  |  |  |  anode-g
*                 |  |  |  |  |  |  |  |  |  | 
.SUBCKT HDSP_H403 1  2  3  4  5  6  7  8  9  10

DA1   7 3 dHDSP_H403
DB1   6 3 dHDSP_H403
DC1   4 3 dHDSP_H403
DD1   2 3 dHDSP_H403
DE1   1 3 dHDSP_H403
DF1   9 3 dHDSP_H403
DG1  10 3 dHDSP_H403
DDP1  5 3 dHDSP_H403

DA2   7 8 dHDSP_H403
DB2   6 8 dHDSP_H403
DC2   4 8 dHDSP_H403
DD2   2 8 dHDSP_H403
DE2   1 8 dHDSP_H403
DF2   9 8 dHDSP_H403
DG2  10 8 dHDSP_H403
DDP2  5 8 dHDSP_H403

.MODEL dHDSP_H403 D
+ (  
+     IS = 3.78006861E-14 
+      N = 2.44553183 
+     RS = 19.51958310 
+     BV = 30
+    IBV = 100u 
+ ) 

.ENDS HDSP_H403
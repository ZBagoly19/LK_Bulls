*  
* Diode Model Produced by Altium Ltd  
* Date:  7-Apr-2004 
*  
* Manufacturer: Agilent  
* Component Name: HDSP-5553  
*  
* Parameters derived from information available in data sheet.  
* 
*                 anode-e
*                 |  anode-d
*                 |  |  common-cathode
*                 |  |  |  anode-c
*                 |  |  |  |  anode-DP
*                 |  |  |  |  |  anode-b
*                 |  |  |  |  |  |  anode-a
*                 |  |  |  |  |  |  |  common-cathode
*                 |  |  |  |  |  |  |  |  anode-f
*                 |  |  |  |  |  |  |  |  |  anode-g
*                 |  |  |  |  |  |  |  |  |  |  
.SUBCKT HDSP_5553 1  2  3  4  5  6  7  8  9  10

DA1   7  3  dHDSP_5553
DB1   6  3  dHDSP_5553
DC1   4  3  dHDSP_5553
DD1   2  3  dHDSP_5553
DE1   1  3  dHDSP_5553
DF1   9  3  dHDSP_5553
DG1  10  3  dHDSP_5553
DDP1  5  3  dHDSP_5553

DA2   7  8  dHDSP_5553
DB2   6  8  dHDSP_5553
DC2   4  8  dHDSP_5553
DD2   2  8  dHDSP_5553
DE2   1  8  dHDSP_5553
DF2   9  8  dHDSP_5553
DG2  10  8  dHDSP_5553
DDP2  5  8  dHDSP_5553

.MODEL dHDSP_5553 D
+ (  
+     IS = 7.07436607E-24 
+      N = 1.24380258 
+     RS = 22.12166762 
+     BV = 30
+    IBV = 100u 
+ )  

.ENDS HDSP_5553
*  
* Diode Model Produced by Altium Ltd  
* Date:  6-Apr-2004 
*  
* Manufacturer: Agilent  
* Component Name: HDSP-5601  
*  
* Parameters derived from information available in data sheet.  
* 
*                 cathode-e
*                 |  cathode-d
*                 |  |  common-anode
*                 |  |  |  cathode-c
*                 |  |  |  |  cathode-DP
*                 |  |  |  |  |  cathode-b
*                 |  |  |  |  |  |  cathode-a
*                 |  |  |  |  |  |  |  common-anode
*                 |  |  |  |  |  |  |  |  cathode-f
*                 |  |  |  |  |  |  |  |  |  cathode-g
*                 |  |  |  |  |  |  |  |  |  | 
.SUBCKT HDSP_5601 1  2  3  4  5  6  7  8  9  10

DA1  3  7 dHDSP_5601
DB1  3  6 dHDSP_5601
DC1  3  4 dHDSP_5601
DD1  3  2 dHDSP_5601
DE1  3  1 dHDSP_5601
DF1  3  9 dHDSP_5601
DG1  3 10 dHDSP_5601
DDP1 3  5 dHDSP_5601

DA2  8  7 dHDSP_5601
DB2  8  6 dHDSP_5601
DC2  8  4 dHDSP_5601
DD2  8  2 dHDSP_5601
DE2  8  1 dHDSP_5601
DF2  8  9 dHDSP_5601
DG2  8 10 dHDSP_5601
DDP2 8  5 dHDSP_5601

.MODEL dHDSP_5601 D
+ (  
+     IS = 1.61114016E-27 
+      N = 1.30291189 
+     RS = 12.83456794 
+     BV = 50 
+    IBV = 100u 
+ )

.ENDS HDSP_5601
*  
* Diode Model Produced by Altium Ltd  
* Date:  3-May-2004 
*  
* Manufacturer: Renesas  
* Component Name: HDSP-A153  
*  
* Parameters derived from information available in data sheet.  
* 
*                 common-cathode
*                 |  anode-f
*                 |  |  anode-g
*                 |  |  |  anode-e
*                 |  |  |  |  anode-d
*                 |  |  |  |  |  common-cathode
*                 |  |  |  |  |  |  anode-DP
*                 |  |  |  |  |  |  |  anode-c
*                 |  |  |  |  |  |  |  |  anode-b
*                 |  |  |  |  |  |  |  |  |  anode-a
*                 |  |  |  |  |  |  |  |  |  |
.SUBCKT HDSP_A153 1  2  3  4  5  6  7  8  9  10

DA1  10  1  dHDSP_A153
DB1   9  1  dHDSP_A153
DC1   8  1  dHDSP_A153
DD1   5  1  dHDSP_A153
DE1   4  1  dHDSP_A153
DF1   2  1  dHDSP_A153
DG1   3  1  dHDSP_A153
DDP1  7  1  dHDSP_A153

DA2  10  6  dHDSP_A153
DB2   9  6  dHDSP_A153
DC2   8  6  dHDSP_A153
DD2   5  6  dHDSP_A153
DE2   4  6  dHDSP_A153
DF2   2  6  dHDSP_A153
DG2   3  6  dHDSP_A153
DDP2  7  6  dHDSP_A153

.MODEL dHDSP_A153 D
+ (  
+    IS  = 2.08276754E-16 
+     N  = 2.17799178 
+    RS  = 0.50892350
+    BV  = 14.25
+   IBV  = 100u
+ )  

.ENDS HDSP_A153
*  
* Diode Model Produced by Altium Ltd  
* Date:  10-Mar-2004 
*  
* Manufacturer: Agilent  
* Component Name: HDSP-303G  
*  
* Parameters derived from information available in data sheet.  
*
*                 anode-G
*                 |  anode-F
*                 |  |  comon-cathode
*                 |  |  |  anode-E
*                 |  |  |  |  anode-D
*                 |  |  |  |  |  anode-DP
*                 |  |  |  |  |  |  anode-C
*                 |  |  |  |  |  |  |  comon-cathode
*                 |  |  |  |  |  |  |  |  anode-B
*                 |  |  |  |  |  |  |  |  |  anode-A
*                 |  |  |  |  |  |  |  |  |  |  
.SUBCKT HDSP_303G 1  2  3  4  5  6  7  8  9  10

DA1  10  3  dHDSP_303G
DB1   9  3  dHDSP_303G
DC1   7  3  dHDSP_303G
DD1   5  3  dHDSP_303G
DE1   4  3  dHDSP_303G
DF1   2  3  dHDSP_303G
DG1   1  3  dHDSP_303G
DDP1  6  3  dHDSP_303G

DA2  10  8  dHDSP_303G
DB2   9  8  dHDSP_303G
DC2   7  8  dHDSP_303G
DD2   5  8  dHDSP_303G
DE2   4  8  dHDSP_303G
DF2   2  8  dHDSP_303G
DG2   1  8  dHDSP_303G
DDP2  6  8  dHDSP_303G

.MODEL dHDSP_303G D
+ (  
+     IS = 3.14401041E-29 
+      N = 1.25233679 
+     RS = 9.99993505 
+     BV = 4.8 
+    IBV = 100u 
+ )  

.ENDS HDSP_303G
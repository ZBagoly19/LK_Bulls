*  
* Diode Model Produced by Altium Ltd  
* Date:  6-Apr-2004 
*  
* Manufacturer: Agilent  
* Component Name: HDSP-5721  
*  
* Parameters derived from information available in data sheet.  
* 
*                 E-cathode-1
*                 |  D-cathode-1
*                 |  |  C-cathode-1
*                 |  |  |  DP-cathode-1
*                 |  |  |  |  E-cathode-1
*                 |  |  |  |  |  D-cathode-2
*                 |  |  |  |  |  |  G-cathode-2
*                 |  |  |  |  |  |  |  C-cathode-2
*                 |  |  |  |  |  |  |  |  DP-cathode-2
*                 |  |  |  |  |  |  |  |  |  B-cathode-2
*                 |  |  |  |  |  |  |  |  |  |  A-cathode-2
*                 |  |  |  |  |  |  |  |  |  |  |  F-cathode-2
*                 |  |  |  |  |  |  |  |  |  |  |  |  common-anode-2
*                 |  |  |  |  |  |  |  |  |  |  |  |  |  common-anode-1
*                 |  |  |  |  |  |  |  |  |  |  |  |  |  |  B-cathode-1
*                 |  |  |  |  |  |  |  |  |  |  |  |  |  |  |  A-cathode-1
*                 |  |  |  |  |  |  |  |  |  |  |  |  |  |  |  |  G-cathode-1
*                 |  |  |  |  |  |  |  |  |  |  |  |  |  |  |  |  |  F-cathode-1
*                 |  |  |  |  |  |  |  |  |  |  |  |  |  |  |  |  |  |
.SUBCKT HDSP_5721 1  2  3  4  5  6  7  8  9  10 11 12 13 14 15 16 17 18

DA1  14  16  dHDSP_5721
DB1  14  15  dHDSP_5721
DC1  14   3  dHDSP_5721
DD1  14   2  dHDSP_5721
DE1  14   1  dHDSP_5721
DF1  14  18  dHDSP_5721
DG1  14  17  dHDSP_5721
DDP1 14   4  dHDSP_5721

DA2  13  11  dHDSP_5721
DB2  13  10  dHDSP_5721
DC2  13   8  dHDSP_5721
DD2  13   6  dHDSP_5721
DE2  13   5  dHDSP_5721
DF2  13  12  dHDSP_5721
DG2  13   7  dHDSP_5721
DDP2 13   9  dHDSP_5721

.MODEL dHDSP_5721 D
+ (  
+     IS = 1.82902372E-24 
+      N = 1.34581490 
+     RS = 23.36447097 
+     BV = 40 
+    IBV = 100u 
+ ) 

.ENDS HDSP_5721
*  
* Diode Model Produced by Altium Ltd  
* Date:  7-Apr-2004 
*  
* Manufacturer: Agilent  
* Component Name: HDSP-516L  
*  
* Parameters derived from information available in data sheet.  
* 
*                 e - anode
*                 |  d - anode
*                 |  |  common-cathode
*                 |  |  |  c - anode
*                 |  |  |  |  DP - anode
*                 |  |  |  |  |  b - anode
*                 |  |  |  |  |  |  a - anode
*                 |  |  |  |  |  |  |  common-cathode
*                 |  |  |  |  |  |  |  |  f - anode
*                 |  |  |  |  |  |  |  |  |  g - anode
*                 |  |  |  |  |  |  |  |  |  | 
.SUBCKT HDSP_516L 1  2  3  4  5  6  7  8  9  10

DA1   7 3 dHDSP_516L
DB1   6 3 dHDSP_516L
DC1   4 3 dHDSP_516L
DD1   2 3 dHDSP_516L
DE1   1 3 dHDSP_516L
DF1   9 3 dHDSP_516L
DG1  10 3 dHDSP_516L
DDP1  5 3 dHDSP_516L

DA2   7 8 dHDSP_516L
DB2   6 8 dHDSP_516L
DC2   4 8 dHDSP_516L
DD2   2 8 dHDSP_516L
DE2   1 8 dHDSP_516L
DF2   9 8 dHDSP_516L
DG2  10 8 dHDSP_516L
DDP2  5 8 dHDSP_516L

.MODEL dHDSP_516L D
+ (  
+     IS = 1.84086967E-50 
+      N = 0.55445364 
+     RS = 251.75
+     BV = 30
+    IBV = 100u 
+ )  

.ENDS HDSP_516L
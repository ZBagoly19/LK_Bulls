*  
* Diode Model Produced by Altium Ltd  
* Date:  10-Mar-2004 
*  
* Manufacturer: Agilent  
* Component Name: HDSP-333Y  
*  
* Parameters derived from information available in data sheet.  
*
*                 anode-F
*                 |  anode-G
*                 |  |  common-cathode
*                 |  |  |  anode-E
*                 |  |  |  |  anode-D
*                 |  |  |  |  |  anode-C
*                 |  |  |  |  |  |  anode-DP
*                 |  |  |  |  |  |  |  common-cathode
*                 |  |  |  |  |  |  |  |  anode-B
*                 |  |  |  |  |  |  |  |  |  anode-A
*                 |  |  |  |  |  |  |  |  |  |  
.SUBCKT HDSP_333Y 1  2  4  6  7  8  9  12 13 14

DA1  14  4  dHDSP_333Y
DB1  13  4  dHDSP_333Y
DC1   8  4  dHDSP_333Y
DD1   7  4  dHDSP_333Y
DE1   6  4  dHDSP_333Y
DF1   1  4  dHDSP_333Y
DG1   2  4  dHDSP_333Y
DDP1  9  4  dHDSP_333Y

DA2  14 12  dHDSP_333Y
DB2  13 12  dHDSP_333Y
DC2   8 12  dHDSP_333Y
DD2   7 12  dHDSP_333Y
DE2   6 12  dHDSP_333Y
DF2   1 12  dHDSP_333Y
DG2   2 12  dHDSP_333Y
DDP2  9 12  dHDSP_333Y

.MODEL dHDSP_333Y D
+ (  
+     IS = 1.56127529E-27 
+      N = 1.25814710 
+     RS = 11.53505957 
+     BV = 4.8 
+    IBV = 100u 
+ )  

.ENDS HDSP_333Y
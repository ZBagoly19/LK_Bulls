*  
* Diode Model Produced by Altium Ltd  
* Date:  7-Apr-2004 
*  
* Manufacturer: Agilent  
* Component Name: HDSP-316Y  
*  
* Parameters derived from information available in data sheet.  
* 
*                 g - anode
*                 |  f - anode
*                 |  |  common-cathode
*                 |  |  |  e - anode
*                 |  |  |  |  d - anode
*                 |  |  |  |  |  DP - anode
*                 |  |  |  |  |  |  c - anode
*                 |  |  |  |  |  |  |  common-cathode
*                 |  |  |  |  |  |  |  |  b - anode
*                 |  |  |  |  |  |  |  |  |  a - anode
*                 |  |  |  |  |  |  |  |  |  | 
.SUBCKT HDSP_316Y 1  2  3  4  5  6  7  8  9  10

DA1  10 3 dHDSP_316Y
DB1   9 3 dHDSP_316Y
DC1   7 3 dHDSP_316Y
DD1   5 3 dHDSP_316Y
DE1   4 3 dHDSP_316Y
DF1   2 3 dHDSP_316Y
DG1   1 3 dHDSP_316Y
DDP1  6 3 dHDSP_316Y

DA2  10 8 dHDSP_316Y
DB2   9 8 dHDSP_316Y
DC2   7 8 dHDSP_316Y
DD2   5 8 dHDSP_316Y
DE2   4 8 dHDSP_316Y
DF2   2 8 dHDSP_316Y
DG2   1 8 dHDSP_316Y
DDP2  6 8 dHDSP_316Y

.MODEL dHDSP_316Y D
+ (  
+     IS = 3.94588412E-15 
+      N = 2.33201916 
+     RS = 23.30053910 
+     BV = 50 
+    IBV = 100u 
+ )  

.ENDS HDSP_316Y
*  
* Diode Model Produced by Altium Ltd  
* Date:  7-Apr-2004 
*  
* Manufacturer: Agilent  
* Component Name: HDSP-316H  
*  
* Parameters derived from information available in data sheet.  
* 
*                 g - anode
*                 |  f - anode
*                 |  |  common-cathode
*                 |  |  |  e - anode
*                 |  |  |  |  d - anode
*                 |  |  |  |  |  DP - anode
*                 |  |  |  |  |  |  c - anode
*                 |  |  |  |  |  |  |  common-cathode
*                 |  |  |  |  |  |  |  |  b - anode
*                 |  |  |  |  |  |  |  |  |  a - anode
*                 |  |  |  |  |  |  |  |  |  | 
.SUBCKT HDSP_316H 1  2  3  4  5  6  7  8  9  10

DA1  10 3 dHDSP_316H
DB1   9 3 dHDSP_316H
DC1   7 3 dHDSP_316H
DD1   5 3 dHDSP_316H
DE1   4 3 dHDSP_316H
DF1   2 3 dHDSP_316H
DG1   1 3 dHDSP_316H
DDP1  6 3 dHDSP_316H

DA2  10 8 dHDSP_316H
DB2   9 8 dHDSP_316H
DC2   7 8 dHDSP_316H
DD2   5 8 dHDSP_316H
DE2   4 8 dHDSP_316H
DF2   2 8 dHDSP_316H
DG2   1 8 dHDSP_316H
DDP2  6 8 dHDSP_316H

.MODEL dHDSP_316H D
+ (  
+    IS  = 2.08276754E-16 
+     N  = 2.17799178 
+    RS  = 0.50892350
+    BV  = 14.25
+   IBV  = 100u
+ )  

.ENDS HDSP_316H
*  
* Diode Model Produced by Altium Ltd  
* Date:  10-Mar-2004 
*  
* Manufacturer: Agilent  
* Component Name: HDSP-U401  
*  
* Parameters derived from information available in data sheet.  
*  
*                  cathode-a 
*                  |  cathode-f 
*                  |  |  cathode-g 
*                  |  |  |  cathode-e 
*                  |  |  |  |  cathode-d 
*                  |  |  |  |  |  cathode-DP 
*                  |  |  |  |  |  |  anode-DP 
*                  |  |  |  |  |  |  |  cathode-c 
*                  |  |  |  |  |  |  |  |  common-anode 
*                  |  |  |  |  |  |  |  |  |  cathode-b
*                  |  |  |  |  |  |  |  |  |  |
.SUBCKT HDSP_U401 1  2  3  4  5  6  7  8  9  10

D1  9  1 dHDSP_U401
D2  9  2 dHDSP_U401
D3  9  3 dHDSP_U401
D4  9  4 dHDSP_U401
D5  9  5 dHDSP_U401
D6  7  6 dHDSP_U401
D7  9  8 dHDSP_U401
D8  9 10 dHDSP_U401

.MODEL dHDSP_U401 D
+ (  
+     IS = 3.04174763E-24 
+      N = 1.23122391 
+     RS = 24.19303791 
+     BV = 30
+    IBV = 100u 
+ )  

.ENDS HDSP_U401
*  
* Diode Model Produced by Altium Ltd  
* Date:  3-May-2004 
*  
* Manufacturer: Renesas  
* Component Name: HDSP-7804  
*  
* Parameters derived from information available in data sheet.  
* 
*                 anode-colon
*                 |  anode-f
*                 |  |  anode-g
*                 |  |  |  anode-e
*                 |  |  |  |  anode-d
*                 |  |  |  |  |  common-cathode
*                 |  |  |  |  |  |  anode-DP
*                 |  |  |  |  |  |  |  anode-c
*                 |  |  |  |  |  |  |  |  anode-b
*                 |  |  |  |  |  |  |  |  |  anode-a
*                 |  |  |  |  |  |  |  |  |  |
.SUBCKT HDSP_7804 1  2  3  4  5  6  7  8  9  10

DA  10  6  dHDSP_7804
DB   9  6  dHDSP_7804
DC   8  6  dHDSP_7804
DD   5  6  dHDSP_7804
DE   4  6  dHDSP_7804
DF   2  6  dHDSP_7804
DG   3  6  dHDSP_7804
DDP  7  6  dHDSP_7804
DCL  1  6  dHDSP_7804

.MODEL dHDSP_7804 D
+ (  
+     IS = 1.61114016E-27 
+      N = 1.30291189 
+     RS = 12.83456794 
+     BV = 50 
+    IBV = 100u 
+ )  

.ENDS HDSP_7804
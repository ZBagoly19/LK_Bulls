*  
* Diode Model Produced by Altium Ltd  
* Date:  10-Mar-2004 
*  
* Manufacturer: Agilent  
* Component Name: HDSP-513G  
*  
* Parameters derived from information available in data sheet.  
*  
*                 anode-e 
*                 |  anode-d 
*                 |  |  common-cathode 
*                 |  |  |  anode-c 
*                 |  |  |  |  anode-DP 
*                 |  |  |  |  |  anode-b 
*                 |  |  |  |  |  |  anode-a 
*                 |  |  |  |  |  |  |  common-cathode 
*                 |  |  |  |  |  |  |  |  anode-f 
*                 |  |  |  |  |  |  |  |  |  anode-g
*                 |  |  |  |  |  |  |  |  |  |
.SUBCKT HDSP_513G 1  2  3  4  5  6  7  8  9  10

DA1  7 3 dHDSP_513G
DB1  6 3 dHDSP_513G
DC1  4 3 dHDSP_513G
DD1  2 3 dHDSP_513G
DE1  1 3 dHDSP_513G
DF1  9 3 dHDSP_513G
DG1 10 3 dHDSP_513G

DA2  7 8 dHDSP_513G
DB2  6 8 dHDSP_513G
DC2  4 8 dHDSP_513G
DD2  2 8 dHDSP_513G
DE2  1 8 dHDSP_513G
DF2  9 8 dHDSP_513G
DG2 10 8 dHDSP_513G

.MODEL dHDSP_513G D
+ (  
+     IS = 1.61114016E-27 
+      N = 1.30291189 
+     RS = 12.83456794 
+     BV = 50 
+    IBV = 100u 
+ )  

.ENDS HDSP_513G
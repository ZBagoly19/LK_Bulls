*  
* Diode Model Produced by Altium Ltd  
* Date:  10-Mar-2004 
*  
* Manufacturer: Agilent  
* Component Name: HDSP-F503  
*  
* Parameters derived from information available in data sheet.  
*  
*                 common-cathode 
*                 |  anode-f 
*                 |  |  anode-g 
*                 |  |  |  anode-e 
*                 |  |  |  |  anode-d 
*                 |  |  |  |  |  common-cathode 
*                 |  |  |  |  |  |  anode-DP 
*                 |  |  |  |  |  |  |  anode-c 
*                 |  |  |  |  |  |  |  |  anode-b 
*                 |  |  |  |  |  |  |  |  |  anode-a
*                 |  |  |  |  |  |  |  |  |  |
.SUBCKT HDSP_F503 1  2  3  4  5  6  7  8  9  10

DA1  10 1 dHDSP_F503
DB1   9 1 dHDSP_F503
DC1   8 1 dHDSP_F503
DD1   5 1 dHDSP_F503
DE1   4 1 dHDSP_F503
DF1   2 1 dHDSP_F503
DG1   3 1 dHDSP_F503
DDP1  7 1 dHDSP_F503

DA2  10 6 dHDSP_F503
DB2   9 6 dHDSP_F503
DC2   8 6 dHDSP_F503
DD2   5 6 dHDSP_F503
DE2   4 6 dHDSP_F503
DF2   2 6 dHDSP_F503
DG2   3 6 dHDSP_F503
DDP2  7 6 dHDSP_F503

.MODEL dHDSP_F503 D
+ (  
+     IS = 1.61114016E-27 
+      N = 1.30291189 
+     RS = 12.83456794 
+     BV = 50 
+    IBV = 100u 
+ ) 

.ENDS HDSP_F503
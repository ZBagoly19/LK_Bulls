*  
* Diode Model Produced by Altium Ltd  
* Date:  10-Mar-2004 
*  
* Manufacturer: Agilent  
* Component Name: HDSP-A111  
*  
* Parameters derived from information available in data sheet.  
*
*                 common-anode
*                 |  cathode-f
*                 |  |  cathode-g
*                 |  |  |  cathode-e
*                 |  |  |  |  cathode-d
*                 |  |  |  |  |  common-anode
*                 |  |  |  |  |  |  cathode-DP
*                 |  |  |  |  |  |  |  cathode-c
*                 |  |  |  |  |  |  |  |  cathode-b
*                 |  |  |  |  |  |  |  |  |  cathode-a
*                 |  |  |  |  |  |  |  |  |  |
.SUBCKT HDSP_A111 1  2  3  4  5  6  7  8  9  10

DA1  1  10 dHDSP_A111
DB1  1   9 dHDSP_A111
DC1  1   8 dHDSP_A111
DD1  1   5 dHDSP_A111
DE1  1   4 dHDSP_A111
DF1  1   2 dHDSP_A111
DG1  1   3 dHDSP_A111
DDP1 1   7 dHDSP_A111

DA2  6  10 dHDSP_A111
DB2  6   9 dHDSP_A111
DC2  6   8 dHDSP_A111
DD2  6   5 dHDSP_A111
DE2  6   4 dHDSP_A111
DF2  6   2 dHDSP_A111
DG2  6   3 dHDSP_A111
DDP2 6   7 dHDSP_A111

.MODEL dHDSP_A111 D
+ (  
+    IS  = 2.08276754E-16 
+     N  = 2.17799178 
+    RS  = 0.50892350
+    BV  = 14.25
+   IBV  = 100u
+ )  

.ENDS HDSP_A111
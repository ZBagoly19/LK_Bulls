*  
* Diode Model Produced by Altium Ltd  
* Date:  7-Apr-2004 
*  
* Manufacturer: Agilent  
* Component Name: HDSP-3600  
*  
* Parameters derived from information available in data sheet.  
* 
*                 cathode-a
*                 |  cathode-f
*                 |  |  common-anode
*                 |  |  |  cathode-DP
*                 |  |  |  |  cathode-e
*                 |  |  |  |  |  cathode-d
*                 |  |  |  |  |  |  cathode-c
*                 |  |  |  |  |  |  |  cathode-g
*                 |  |  |  |  |  |  |  |  cathode-b
*                 |  |  |  |  |  |  |  |  |  common-anode
*                 |  |  |  |  |  |  |  |  |  |
*                 |  |  |  |  |  |  |  |  |  | 
.SUBCKT HDSP_3600 1  2  3  6  7  8  10 11 13 14

DA1   3  1 dHDSP_3600
DB1   3 13 dHDSP_3600
DC1   3 10 dHDSP_3600
DD1   3  8 dHDSP_3600
DE1   3  7 dHDSP_3600
DF1   3  2 dHDSP_3600
DG1   3 11 dHDSP_3600
DDP1  3  6 dHDSP_3600

DA2  14  1 dHDSP_3600
DB2  14 13 dHDSP_3600
DC2  14 10 dHDSP_3600
DD2  14  8 dHDSP_3600
DE2  14  7 dHDSP_3600
DF2  14  2 dHDSP_3600
DG2  14 11 dHDSP_3600
DDP2 14  6 dHDSP_3600


.MODEL dHDSP_3600 D
+ (  
+     IS = 1.61114016E-27 
+      N = 1.30291189 
+     RS = 12.83456794 
+     BV = 50 
+    IBV = 100u 
+ )  

.ENDS HDSP_3600
*  
* Diode Model Produced by Altium Ltd  
* Date:  3-May-2004 
*  
* Manufacturer: Renesas  
* Component Name: HDSP-A151  
*  
* Parameters derived from information available in data sheet.  
* 
*                 common-anode
*                 |  cathode-f
*                 |  |  cathode-g
*                 |  |  |  cathode-e
*                 |  |  |  |  cathode-d
*                 |  |  |  |  |  common-anode
*                 |  |  |  |  |  |  cathode-DP
*                 |  |  |  |  |  |  |  cathode-c
*                 |  |  |  |  |  |  |  |  cathode-b
*                 |  |  |  |  |  |  |  |  |  cathode-a
*                 |  |  |  |  |  |  |  |  |  |
.SUBCKT HDSP_A151 1  2  3  4  5  6  7  8  9  10

DA1  1  10  dHDSP_A151
DB1  1   9  dHDSP_A151
DC1  1   8  dHDSP_A151
DD1  1   5  dHDSP_A151
DE1  1   4  dHDSP_A151
DF1  1   2  dHDSP_A151
DG1  1   3  dHDSP_A151
DDP1 1   7  dHDSP_A151

DA2  6  10  dHDSP_A151
DB2  6   9  dHDSP_A151
DC2  6   8  dHDSP_A151
DD2  6   5  dHDSP_A151
DE2  6   4  dHDSP_A151
DF2  6   2  dHDSP_A151
DG2  6   3  dHDSP_A151
DDP2 6   7  dHDSP_A151

.MODEL dHDSP_A151 D
+ (  
+    IS  = 2.08276754E-16 
+     N  = 2.17799178 
+    RS  = 0.50892350
+    BV  = 14.25
+   IBV  = 100u
+ )  

.ENDS HDSP_A151
*  
* Diode Model Produced by Altium Ltd  
* Date:  7-Apr-2004 
*  
* Manufacturer: Agilent  
* Component Name: HDSP-315E  
*  
* Parameters derived from information available in data sheet.  
* 
*                 g - cathode
*                 |  f - cathode
*                 |  |  common-anode
*                 |  |  |  e - cathode
*                 |  |  |  |  d - cathode
*                 |  |  |  |  |  DP - cathode
*                 |  |  |  |  |  |  c - cathode
*                 |  |  |  |  |  |  |  common-anode
*                 |  |  |  |  |  |  |  |  b - cathode
*                 |  |  |  |  |  |  |  |  |  a - cathode
*                 |  |  |  |  |  |  |  |  |  | 
.SUBCKT HDSP_315E 1  2  3  4  5  6  7  8  9  10

DA1  3 10 dHDSP_315E
DB1  3  9 dHDSP_315E
DC1  3  7 dHDSP_315E
DD1  3  5 dHDSP_315E
DE1  3  4 dHDSP_315E
DF1  3  2 dHDSP_315E
DG1  3  1 dHDSP_315E
DDP1 3  6 dHDSP_315E

DA2  8 10 dHDSP_315E
DB2  8  9 dHDSP_315E
DC2  8  7 dHDSP_315E
DD2  8  5 dHDSP_315E
DE2  8  4 dHDSP_315E
DF2  8  2 dHDSP_315E
DG2  8  1 dHDSP_315E
DDP2 8  6 dHDSP_315E

.MODEL dHDSP_315E D
+ (  
+     IS = 1.21481726E-49 
+      N = 0.55445364 
+     RS = 25.38287000 
+     BV = 30
+    IBV = 100u 
+ )  

.ENDS HDSP_315E
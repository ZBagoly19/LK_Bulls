*  
* Diode Model Produced by Altium Ltd  
* Date:  10-Mar-2004 
*  
* Manufacturer: Agilent  
* Component Name: HDSP-313Y  
*  
* Parameters derived from information available in data sheet.  
*  
*                 anode-G 
*                 |  anode-F 
*                 |  |  common-cathode 
*                 |  |  |  anode-E 
*                 |  |  |  |  anode-D 
*                 |  |  |  |  |  anode-DP 
*                 |  |  |  |  |  |  anode-C 
*                 |  |  |  |  |  |  |  common-cathode 
*                 |  |  |  |  |  |  |  |  anode-B 
*                 |  |  |  |  |  |  |  |  |  anode-A
*                 |  |  |  |  |  |  |  |  |  |
.SUBCKT HDSP_313Y 1  2  3  4  5  6  7  8  9  10

DA1  3  10 dHDSP_313Y
DB1  3   9 dHDSP_313Y
DC1  3   7 dHDSP_313Y
DD1  3   5 dHDSP_313Y
DE1  3   4 dHDSP_313Y
DF1  3   2 dHDSP_313Y
DG1  3   1 dHDSP_313Y
DDP1 3   6 dHDSP_313Y

DA2  8  10 dHDSP_313Y
DB2  8   9 dHDSP_313Y
DC2  8   7 dHDSP_313Y
DD2  8   5 dHDSP_313Y
DE2  8   4 dHDSP_313Y
DF2  8   2 dHDSP_313Y
DG2  8   1 dHDSP_313Y
DDP2 8   6 dHDSP_313Y

.MODEL dHDSP_313Y D
+ (  
+     IS = 1.56127529E-27 
+      N = 1.25814710 
+     RS = 11.53505957 
+     BV = 4.8 
+    IBV = 100u 
+ )   

.ENDS HDSP_313Y
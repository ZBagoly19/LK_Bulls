*  
* Diode Model Produced by Altium Ltd  
* Date:  3-May-2004 
*  
* Manufacturer: Renesas  
* Component Name: HDSP-7802  
*  
* Parameters derived from information available in data sheet.  
* 
*                 cathode-colon
*                 |  cathode-f
*                 |  |  cathode-g
*                 |  |  |  cathode-e
*                 |  |  |  |  cathode-d
*                 |  |  |  |  |  common-anode
*                 |  |  |  |  |  |  cathode-DP
*                 |  |  |  |  |  |  |  cathode-c
*                 |  |  |  |  |  |  |  |  cathode-b
*                 |  |  |  |  |  |  |  |  |  cathode-a
*                 |  |  |  |  |  |  |  |  |  |
.SUBCKT HDSP_7802 1  2  3  4  5  6  7  8  9  10

DA  6  10  dHDSP_7802
DB  6   9  dHDSP_7802
DC  6   8  dHDSP_7802
DD  6   5  dHDSP_7802
DE  6   4  dHDSP_7802
DF  6   2  dHDSP_7802
DG  6   3  dHDSP_7802
DDP 6   7  dHDSP_7802
DCL 6   1  dHDSP_7802

.MODEL dHDSP_7802 D
+ (  
+     IS = 1.61114016E-27 
+      N = 1.30291189 
+     RS = 12.83456794 
+     BV = 50 
+    IBV = 100u 
+ )  

.ENDS HDSP_7802
*  
* Diode Model Produced by Altium Ltd  
* Date:  7-Apr-2004 
*  
* Manufacturer: Agilent  
* Component Name: HDSP-4205  
*  
* Parameters derived from information available in data sheet.  
* 
*                 anode-a 
*                 |  anode-f 
*                 |  |  common-cathode
*                 |  |  |  anode-e 
*                 |  |  |  |  common-cathode 
*                 |  |  |  |  |  anode-DP 
*                 |  |  |  |  |  |  anode-d 
*                 |  |  |  |  |  |  |  common-cathode 
*                 |  |  |  |  |  |  |  |  anode-c 
*                 |  |  |  |  |  |  |  |  |  anode-g 
*                 |  |  |  |  |  |  |  |  |  |  anode-b 
*                 |  |  |  |  |  |  |  |  |  |  |  common-cathode
*                 |  |  |  |  |  |  |  |  |  |  |  |
.SUBCKT HDSP_4205 2  3  4  5  6  7  11 12 13 14 15 17

DA1   2  4 dHDSP_4205
DB1  15  4 dHDSP_4205
DC1  13  4 dHDSP_4205
DD1  11  4 dHDSP_4205
DE1   5  4 dHDSP_4205
DF1   3  4 dHDSP_4205
DG1  14  4 dHDSP_4205
DDP1  7  4 dHDSP_4205

DA2   2  6 dHDSP_4205
DB2  15  6 dHDSP_4205
DC2  13  6 dHDSP_4205
DD2  11  6 dHDSP_4205
DE2   5  6 dHDSP_4205
DF2   3  6 dHDSP_4205
DG2  14  6 dHDSP_4205
DDP2  7  6 dHDSP_4205

DA3   2 12 dHDSP_4205
DB3  15 12 dHDSP_4205
DC3  13 12 dHDSP_4205
DD3  11 12 dHDSP_4205
DE3   5 12 dHDSP_4205
DF3   3 12 dHDSP_4205
DG3  14 12 dHDSP_4205
DDP3  7 12 dHDSP_4205

DA4   2 17 dHDSP_4205
DB4  15 17 dHDSP_4205
DC4  13 17 dHDSP_4205
DD4  11 17 dHDSP_4205
DE4   5 17 dHDSP_4205
DF4   3 17 dHDSP_4205
DG4  14 17 dHDSP_4205
DDP4  7 17 dHDSP_4205


.MODEL dHDSP_4205 D
+ (  
+     IS = 8.07922028E-13 
+      N = 3.08151986 
+     RS = 5.65168121 
+     BV = 2.25
+    IBV = 100u 
+ )  

.ENDS HDSP_4205
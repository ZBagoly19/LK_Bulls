*  
* Diode Model Produced by Altium Ltd  
* Date:  7-Apr-2004 
*  
* Manufacturer: Agilent  
* Component Name: HDSP-4200  
*  
* Parameters derived from information available in data sheet.  
* 
*                 cathode-a 
*                 |  cathode-f 
*                 |  |  common-anode
*                 |  |  |  cathode-e 
*                 |  |  |  |  common-anode 
*                 |  |  |  |  |  cathode-DP 
*                 |  |  |  |  |  |  cathode-d 
*                 |  |  |  |  |  |  |  common-anode 
*                 |  |  |  |  |  |  |  |  cathode-c 
*                 |  |  |  |  |  |  |  |  |  cathode-g 
*                 |  |  |  |  |  |  |  |  |  |  cathode-b 
*                 |  |  |  |  |  |  |  |  |  |  |  common-anode
*                 |  |  |  |  |  |  |  |  |  |  |  |
.SUBCKT HDSP_4200 2  3  4  5  6  7  11 12 13 14 15 17

DA1   4  2 dHDSP_4200
DB1   4 15 dHDSP_4200
DC1   4 13 dHDSP_4200
DD1   4 11 dHDSP_4200
DE1   4  5 dHDSP_4200
DF1   4  3 dHDSP_4200
DG1   4 14 dHDSP_4200
DDP1  4  7 dHDSP_4200

DA2   6  2 dHDSP_4200
DB2   6 15 dHDSP_4200
DC2   6 13 dHDSP_4200
DD2   6 11 dHDSP_4200
DE2   6  5 dHDSP_4200
DF2   6  3 dHDSP_4200
DG2   6 14 dHDSP_4200
DDP2  6  7 dHDSP_4200

DA3  12  2 dHDSP_4200
DB3  12 15 dHDSP_4200
DC3  12 13 dHDSP_4200
DD3  12 11 dHDSP_4200
DE3  12  5 dHDSP_4200
DF3  12  3 dHDSP_4200
DG3  12 14 dHDSP_4200
DDP3 12  7 dHDSP_4200

DA4  17  2 dHDSP_4200
DB4  17 15 dHDSP_4200
DC4  17 13 dHDSP_4200
DD4  17 11 dHDSP_4200
DE4  17  5 dHDSP_4200
DF4  17  3 dHDSP_4200
DG4  17 14 dHDSP_4200
DDP4 17  7 dHDSP_4200


.MODEL dHDSP_4200 D
+ (  
+     IS = 8.07922028E-13 
+      N = 3.08151986 
+     RS = 5.65168121 
+     BV = 2.25
+    IBV = 100u 
+ )  

.ENDS HDSP_4200
*  
* Diode Model Produced by Altium Ltd  
* Date:  10-Mar-2004 
*  
* Manufacturer: Agilent  
* Component Name: HDSP-F203  
*  
* Parameters derived from information available in data sheet.  
*  
*                 common-cathode 
*                 |  anode-f 
*                 |  |  anode-g 
*                 |  |  |  anode-e 
*                 |  |  |  |  anode-d 
*                 |  |  |  |  |  common-cathode 
*                 |  |  |  |  |  |  anode-DP 
*                 |  |  |  |  |  |  |  anode-c 
*                 |  |  |  |  |  |  |  |  anode-b 
*                 |  |  |  |  |  |  |  |  |  anode-a
*                 |  |  |  |  |  |  |  |  |  |
.SUBCKT HDSP_F203 1  2  3  4  5  6  7  8  9  10

DA1  10 1 dHDSP_F203
DB1   9 1 dHDSP_F203
DC1   8 1 dHDSP_F203
DD1   5 1 dHDSP_F203
DE1   4 1 dHDSP_F203
DF1   2 1 dHDSP_F203
DG1   3 1 dHDSP_F203
DDP1  7 1 dHDSP_F203

DA2  10 6 dHDSP_F203
DB2   9 6 dHDSP_F203
DC2   8 6 dHDSP_F203
DD2   5 6 dHDSP_F203
DE2   4 6 dHDSP_F203
DF2   2 6 dHDSP_F203
DG2   3 6 dHDSP_F203
DDP2  7 6 dHDSP_F203

.MODEL dHDSP_F203 D
+ (  
+     IS = 3.04174763E-24 
+      N = 1.23122391 
+     RS = 24.19303791 
+     BV = 30
+    IBV = 100u 
+ )  

.ENDS HDSP_F203
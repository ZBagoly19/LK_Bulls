*  
* Diode Model Produced by Altium Ltd  
* Date:  10-Mar-2004 
*  
* Manufacturer: Agilent  
* Component Name: HDSP-513Y  
*  
* Parameters derived from information available in data sheet.  
*  
*                 anode-e 
*                 |  anode-d 
*                 |  |  common-cathode 
*                 |  |  |  anode-c 
*                 |  |  |  |  anode-DP 
*                 |  |  |  |  |  anode-b 
*                 |  |  |  |  |  |  anode-a 
*                 |  |  |  |  |  |  |  common-cathode 
*                 |  |  |  |  |  |  |  |  anode-f 
*                 |  |  |  |  |  |  |  |  |  anode-g
*                 |  |  |  |  |  |  |  |  |  |
.SUBCKT HDSP_513Y 1  2  3  4  5  6  7  8  9  10

DA1  7 3 dHDSP_513Y
DB1  6 3 dHDSP_513Y
DC1  4 3 dHDSP_513Y
DD1  2 3 dHDSP_513Y
DE1  1 3 dHDSP_513Y
DF1  9 3 dHDSP_513Y
DG1 10 3 dHDSP_513Y

DA2  7 8 dHDSP_513Y
DB2  6 8 dHDSP_513Y
DC2  4 8 dHDSP_513Y
DD2  2 8 dHDSP_513Y
DE2  1 8 dHDSP_513Y
DF2  9 8 dHDSP_513Y
DG2 10 8 dHDSP_513Y

.MODEL dHDSP_513Y D
+ (  
+     IS = 1.56127529E-27 
+      N = 1.25814710 
+     RS = 11.53505957 
+     BV = 4.8 
+    IBV = 100u 
+ )  

.ENDS HDSP_513Y
*  
* Diode Model Produced by Altium Ltd  
* Date:  6-Apr-2004 
*  
* Manufacturer: Agilent  
* Component Name: HDSP-5503  
*  
* Parameters derived from information available in data sheet.  
* 
*                 anode-e
*                 |  anode-d
*                 |  |  common-cathode
*                 |  |  |  anode-c
*                 |  |  |  |  anode-DP
*                 |  |  |  |  |  anode-b
*                 |  |  |  |  |  |  anode-a
*                 |  |  |  |  |  |  |  common-cathode
*                 |  |  |  |  |  |  |  |  anode-f
*                 |  |  |  |  |  |  |  |  |  anode-g
*                 |  |  |  |  |  |  |  |  |  | 
.SUBCKT HDSP_5503 1  2  3  4  5  6  7  8  9  10

DA1   7 3 dHDSP_5503
DB1   6 3 dHDSP_5503
DC1   4 3 dHDSP_5503
DD1   2 3 dHDSP_5503
DE1   1 3 dHDSP_5503
DF1   9 3 dHDSP_5503
DG1  10 3 dHDSP_5503
DDP1  5 3 dHDSP_5503

DA2   7 8 dHDSP_5503
DB2   6 8 dHDSP_5503
DC2   4 8 dHDSP_5503
DD2   2 8 dHDSP_5503
DE2   1 8 dHDSP_5503
DF2   9 8 dHDSP_5503
DG2  10 8 dHDSP_5503
DDP2  5 8 dHDSP_5503

.MODEL dHDSP_5503 D
+ (  
+     IS = 3.78006861E-14 
+      N = 2.44553183 
+     RS = 19.51958310 
+     BV = 30
+    IBV = 100u 
+ )  

.ENDS HDSP_5503
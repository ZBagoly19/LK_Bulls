*  
* Diode Model Produced by Altium Ltd  
* Date:  10-Mar-2004 
*  
* Manufacturer: Agilent  
* Component Name: HDSP-563A  
*  
* Parameters derived from information available in data sheet.  
*
*                 anode-E
*                 |  anode-D
*                 |  |  comon-cathode
*                 |  |  |  anode-C
*                 |  |  |  |  anode-DP
*                 |  |  |  |  |  anode-B
*                 |  |  |  |  |  |  anode-A
*                 |  |  |  |  |  |  |  comon-cathode
*                 |  |  |  |  |  |  |  |  anode-F
*                 |  |  |  |  |  |  |  |  |  anode-G
*                 |  |  |  |  |  |  |  |  |  |  
.SUBCKT HDSP_563A 1  2  3  4  5  6  7  8  9  10

DA1   7  3  dHDSP_563A
DB1   6  3  dHDSP_563A
DC1   4  3  dHDSP_563A
DD1   2  3  dHDSP_563A
DE1   1  3  dHDSP_563A
DF1   9  3  dHDSP_563A
DG1  10  3  dHDSP_563A
DDP1  5  3  dHDSP_563A

DA2   7  8  dHDSP_563A
DB2   6  8  dHDSP_563A
DC2   4  8  dHDSP_563A
DD2   2  8  dHDSP_563A
DE2   1  8  dHDSP_563A
DF2   9  8  dHDSP_563A
DG2  10  8  dHDSP_563A
DDP2  5  8  dHDSP_563A

.MODEL dHDSP_563A D
+ (  
+    IS = 4.59961571E-15 
+     N = 2.40621673 
+    RS = 1.90931135 
+    BV = 4.5
+   IBV = 100u
+ )  

.ENDS HDSP_563A
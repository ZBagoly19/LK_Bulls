*  
* Diode Model Produced by Altium Ltd  
* Date:  7-Apr-2004 
*  
* Manufacturer: Agilent  
* Component Name: HDSP-7511  
*  
* Parameters derived from information available in data sheet.  
*  
*                 common-anode
*                 |  cathode-f
*                 |  |  cathode-g
*                 |  |  |  cathode-e
*                 |  |  |  |  cathode-d
*                 |  |  |  |  |  common-anode
*                 |  |  |  |  |  |  cathode-DP
*                 |  |  |  |  |  |  |  cathode-c
*                 |  |  |  |  |  |  |  |  cathode-b
*                 |  |  |  |  |  |  |  |  |  cathode-a
*                 |  |  |  |  |  |  |  |  |  |
.SUBCKT HDSP_7511 1  2  3  4  5  6  7  8  9  10

DA1  1  10 dHDSP_7511
DB1  1   9 dHDSP_7511
DC1  1   8 dHDSP_7511
DD1  1   5 dHDSP_7511
DE1  1   4 dHDSP_7511
DF1  1   2 dHDSP_7511
DG1  1   3 dHDSP_7511
DDP1 1   7 dHDSP_7511

DA2  6  10 dHDSP_7511
DB2  6   9 dHDSP_7511
DC2  6   8 dHDSP_7511
DD2  6   5 dHDSP_7511
DE2  6   4 dHDSP_7511
DF2  6   2 dHDSP_7511
DG2  6   3 dHDSP_7511
DDP2 6   7 dHDSP_7511

.MODEL dHDSP_7511 D
+ (  
+     IS = 7.07436607E-24 
+      N = 1.24380258 
+     RS = 22.12166762 
+     BV = 30
+    IBV = 100u 
+ )  

.ENDS HDSP_7511
*  
* Diode Model Produced by Altium Ltd  
* Date:  10-Mar-2004 
*  
* Manufacturer: Agilent  
* Component Name: HDSP-H511  
*  
* Parameters derived from information available in data sheet.  
* 
*                 cathode-e
*                 |  cathode-d
*                 |  |  common-anode
*                 |  |  |  cathode-c
*                 |  |  |  |  cathode-DP
*                 |  |  |  |  |  cathode-b
*                 |  |  |  |  |  |  cathode-a
*                 |  |  |  |  |  |  |  common-anode
*                 |  |  |  |  |  |  |  |  cathode-f
*                 |  |  |  |  |  |  |  |  |  cathode-g
*                 |  |  |  |  |  |  |  |  |  | 
.SUBCKT HDSP_H511 1  2  3  4  5  6  7  8  9  10

DA1   3  7  dHDSP_H511
DB1   3  6  dHDSP_H511
DC1   3  4  dHDSP_H511
DD1   3  2  dHDSP_H511
DE1   3  1  dHDSP_H511
DF1   3  9  dHDSP_H511
DG1   3 10  dHDSP_H511
DDP1  3  5  dHDSP_H511

DA2   8  7  dHDSP_H511
DB2   8  6  dHDSP_H511
DC2   8  4  dHDSP_H511
DD2   8  2  dHDSP_H511
DE2   8  1  dHDSP_H511
DF2   8  9  dHDSP_H511
DG2   8 10  dHDSP_H511
DDP2  8  5  dHDSP_H511

.MODEL dHDSP_H511 D
+ (  
+     IS = 1.61114016E-27 
+      N = 1.30291189 
+     RS = 12.83456794 
+     BV = 50 
+    IBV = 100u 
+ )  

.ENDS HDSP_H511
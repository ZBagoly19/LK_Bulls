*  
* Diode Model Produced by Altium Ltd  
* Date:  7-Apr-2004 
*  
* Manufacturer: Agilent  
* Component Name: HDSP-3900  
*  
* Parameters derived from information available in data sheet.  
* 
*                 cathode-a 
*                 |  cathode-f 
*                 |  |  common-anode
*                 |  |  |  cathode-e 
*                 |  |  |  |  common-anode 
*                 |  |  |  |  |  cathode-DP 
*                 |  |  |  |  |  |  cathode-d 
*                 |  |  |  |  |  |  |  common-anode 
*                 |  |  |  |  |  |  |  |  cathode-c 
*                 |  |  |  |  |  |  |  |  |  cathode-g 
*                 |  |  |  |  |  |  |  |  |  |  cathode-b 
*                 |  |  |  |  |  |  |  |  |  |  |  common-anode
*                 |  |  |  |  |  |  |  |  |  |  |  |
.SUBCKT HDSP_3900 2  3  4  5  6  7  11 12 13 14 15 17

DA1   4  2 dHDSP_3900
DB1   4 15 dHDSP_3900
DC1   4 13 dHDSP_3900
DD1   4 11 dHDSP_3900
DE1   4  5 dHDSP_3900
DF1   4  3 dHDSP_3900
DG1   4 14 dHDSP_3900
DDP1  4  7 dHDSP_3900

DA2   6  2 dHDSP_3900
DB2   6 15 dHDSP_3900
DC2   6 13 dHDSP_3900
DD2   6 11 dHDSP_3900
DE2   6  5 dHDSP_3900
DF2   6  3 dHDSP_3900
DG2   6 14 dHDSP_3900
DDP2  6  7 dHDSP_3900

DA3  12  2 dHDSP_3900
DB3  12 15 dHDSP_3900
DC3  12 13 dHDSP_3900
DD3  12 11 dHDSP_3900
DE3  12  5 dHDSP_3900
DF3  12  3 dHDSP_3900
DG3  12 14 dHDSP_3900
DDP3 12  7 dHDSP_3900

DA4  17  2 dHDSP_3900
DB4  17 15 dHDSP_3900
DC4  17 13 dHDSP_3900
DD4  17 11 dHDSP_3900
DE4  17  5 dHDSP_3900
DF4  17  3 dHDSP_3900
DG4  17 14 dHDSP_3900
DDP4 17  7 dHDSP_3900


.MODEL dHDSP_3900 D
+ (  
+     IS = 1E-13 
+      N = 2.7
+     RS = 6.22331865 
+     BV = 2.25
+    IBV = 100u 
+ )  

.ENDS HDSP_3900
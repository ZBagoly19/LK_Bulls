*  
* Diode Model Produced by Altium Ltd  
* Date:  7-Apr-2004 
*  
* Manufacturer: Agilent  
* Component Name: HDSP-516G  
*  
* Parameters derived from information available in data sheet.  
* 
*                 e - anode
*                 |  d - anode
*                 |  |  common-cathode
*                 |  |  |  c - anode
*                 |  |  |  |  DP - anode
*                 |  |  |  |  |  b - anode
*                 |  |  |  |  |  |  a - anode
*                 |  |  |  |  |  |  |  common-cathode
*                 |  |  |  |  |  |  |  |  f - anode
*                 |  |  |  |  |  |  |  |  |  g - anode
*                 |  |  |  |  |  |  |  |  |  | 
.SUBCKT HDSP_516G 1  2  3  4  5  6  7  8  9  10

DA1   7 3 dHDSP_516G
DB1   6 3 dHDSP_516G
DC1   4 3 dHDSP_516G
DD1   2 3 dHDSP_516G
DE1   1 3 dHDSP_516G
DF1   9 3 dHDSP_516G
DG1  10 3 dHDSP_516G
DDP1  5 3 dHDSP_516G

DA2   7 8 dHDSP_516G
DB2   6 8 dHDSP_516G
DC2   4 8 dHDSP_516G
DD2   2 8 dHDSP_516G
DE2   1 8 dHDSP_516G
DF2   9 8 dHDSP_516G
DG2  10 8 dHDSP_516G
DDP2  5 8 dHDSP_516G

.MODEL dHDSP_516G D
+ (  
+     IS = 1.61114016E-27 
+      N = 1.30291189 
+     RS = 12.83456794 
+     BV = 50 
+    IBV = 100u 
+ )  

.ENDS HDSP_516G
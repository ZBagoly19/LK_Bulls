*  
* Diode Model Produced by Altium Ltd  
* Date:  7-Apr-2004 
*  
* Manufacturer: Agilent  
* Component Name: HDSP-515L  
*  
* Parameters derived from information available in data sheet.  
* 
*                 e - cathode
*                 |  d - cathode
*                 |  |  common-anode
*                 |  |  |  c - cathode
*                 |  |  |  |  DP - cathode
*                 |  |  |  |  |  b - cathode
*                 |  |  |  |  |  |  a - cathode
*                 |  |  |  |  |  |  |  common-anode
*                 |  |  |  |  |  |  |  |  f - cathode
*                 |  |  |  |  |  |  |  |  |  g - cathode
*                 |  |  |  |  |  |  |  |  |  | 
.SUBCKT HDSP_515L 1  2  3  4  5  6  7  8  9  10

DA1  3  7 dHDSP_515L
DB1  3  6 dHDSP_515L
DC1  3  4 dHDSP_515L
DD1  3  2 dHDSP_515L
DE1  3  1 dHDSP_515L
DF1  3  9 dHDSP_515L
DG1  3 10 dHDSP_515L
DDP1 3  5 dHDSP_515L

DA2  8  7 dHDSP_515L
DB2  8  6 dHDSP_515L
DC2  8  4 dHDSP_515L
DD2  8  2 dHDSP_515L
DE2  8  1 dHDSP_515L
DF2  8  9 dHDSP_515L
DG2  8 10 dHDSP_515L
DDP2 8  5 dHDSP_515L

.MODEL dHDSP_515L D
+ (  
+     IS = 1.84086967E-50 
+      N = 0.55445364 
+     RS = 251.75
+     BV = 30
+    IBV = 100u 
+ )  

.ENDS HDSP_515L
*  
* Diode Model Produced by Altium Ltd  
* Date:  10-Mar-2004 
*  
* Manufacturer: Agilent  
* Component Name: HDSP-303E  
*  
* Parameters derived from information available in data sheet.  
*
*                 anode-G
*                 |  anode-F
*                 |  |  comon-cathode
*                 |  |  |  anode-E
*                 |  |  |  |  anode-D
*                 |  |  |  |  |  anode-DP
*                 |  |  |  |  |  |  anode-C
*                 |  |  |  |  |  |  |  comon-cathode
*                 |  |  |  |  |  |  |  |  anode-B
*                 |  |  |  |  |  |  |  |  |  anode-A
*                 |  |  |  |  |  |  |  |  |  |  
.SUBCKT HDSP_303E 1  2  3  4  5  6  7  8  9  10

DA1  10  3  dHDSP_303E
DB1   9  3  dHDSP_303E
DC1   7  3  dHDSP_303E
DD1   5  3  dHDSP_303E
DE1   4  3  dHDSP_303E
DF1   2  3  dHDSP_303E
DG1   1  3  dHDSP_303E
DDP1  6  3  dHDSP_303E

DA2  10  8  dHDSP_303E
DB2   9  8  dHDSP_303E
DC2   7  8  dHDSP_303E
DD2   5  8  dHDSP_303E
DE2   4  8  dHDSP_303E
DF2   2  8  dHDSP_303E
DG2   1  8  dHDSP_303E
DDP2  6  8  dHDSP_303E

.MODEL dHDSP_303E D
+ (  
+     IS = 1.37607512E-24 
+      N = 1.38335616 
+     RS = 6.06238569 
+     BV = 4.8 
+    IBV = 100u 
+ ) 

.ENDS HDSP_303E
*  
* Diode Model Produced by Altium Ltd  
* Date:  10-Mar-2004 
*  
* Manufacturer: Agilent  
* Component Name: HDSP-F303  
*  
* Parameters derived from information available in data sheet.  
*  
*                 common-cathode 
*                 |  anode-f 
*                 |  |  anode-g 
*                 |  |  |  anode-e 
*                 |  |  |  |  anode-d 
*                 |  |  |  |  |  common-cathode 
*                 |  |  |  |  |  |  anode-DP 
*                 |  |  |  |  |  |  |  anode-c 
*                 |  |  |  |  |  |  |  |  anode-b 
*                 |  |  |  |  |  |  |  |  |  anode-a
*                 |  |  |  |  |  |  |  |  |  |
.SUBCKT HDSP_F303 1  2  3  4  5  6  7  8  9  10

DA1  10 1 dHDSP_F303
DB1   9 1 dHDSP_F303
DC1   8 1 dHDSP_F303
DD1   5 1 dHDSP_F303
DE1   4 1 dHDSP_F303
DF1   2 1 dHDSP_F303
DG1   3 1 dHDSP_F303
DDP1  7 1 dHDSP_F303

DA2  10 6 dHDSP_F303
DB2   9 6 dHDSP_F303
DC2   8 6 dHDSP_F303
DD2   5 6 dHDSP_F303
DE2   4 6 dHDSP_F303
DF2   2 6 dHDSP_F303
DG2   3 6 dHDSP_F303
DDP2  7 6 dHDSP_F303

.MODEL dHDSP_F303 D
+ (  
+     IS = 6.04055825E-18 
+      N = 1.90788337 
+     RS = 23.52447762 
+     BV = 40
+    IBV = 100u 
+ )  

.ENDS HDSP_F303
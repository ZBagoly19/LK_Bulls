*  
* Diode Model Produced by Altium Ltd  
* Date:  7-Apr-2004 
*  
* Manufacturer: Agilent  
* Component Name: HDSP-A801  
*  
* Parameters derived from information available in data sheet.  
*  
*                 common-anode
*                 |  cathode-f
*                 |  |  cathode-g
*                 |  |  |  cathode-e
*                 |  |  |  |  cathode-d
*                 |  |  |  |  |  common-anode
*                 |  |  |  |  |  |  cathode-DP
*                 |  |  |  |  |  |  |  cathode-c
*                 |  |  |  |  |  |  |  |  cathode-b
*                 |  |  |  |  |  |  |  |  |  cathode-a
*                 |  |  |  |  |  |  |  |  |  |
.SUBCKT HDSP_A801 1  2  3  4  5  6  7  8  9  10

DA1  1  10 dHDSP_A801
DB1  1   9 dHDSP_A801
DC1  1   8 dHDSP_A801
DD1  1   5 dHDSP_A801
DE1  1   4 dHDSP_A801
DF1  1   2 dHDSP_A801
DG1  1   3 dHDSP_A801
DDP1 1   7 dHDSP_A801

DA2  6  10 dHDSP_A801
DB2  6   9 dHDSP_A801
DC2  6   8 dHDSP_A801
DD2  6   5 dHDSP_A801
DE2  6   4 dHDSP_A801
DF2  6   2 dHDSP_A801
DG2  6   3 dHDSP_A801
DDP2 6   7 dHDSP_A801

.MODEL dHDSP_A801 D
+ (  
+     IS = 6.64511693E-21 
+      N = 1.66825537 
+     RS = 20.13814139 
+     BV = 30
+    IBV = 100u 
+ )  

.ENDS HDSP_A801
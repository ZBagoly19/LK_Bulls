*  
* Diode Model Produced by Altium Ltd  
* Date:  7-Apr-2004 
*  
* Manufacturer: Agilent  
* Component Name: HDSP-8600  
*  
* Parameters derived from information available in data sheet.  
*  
*                 cathode-a 
*                 |  cathode-f 
*                 |  |  common-anode 
*                 |  |  |  cathode-e 
*                 |  |  |  |  common-anode 
*                 |  |  |  |  |  cathode-DP 
*                 |  |  |  |  |  |  cathode-d 
*                 |  |  |  |  |  |  |  common-anode 
*                 |  |  |  |  |  |  |  |  cathode-c 
*                 |  |  |  |  |  |  |  |  |  cathode-g 
*                 |  |  |  |  |  |  |  |  |  |  cathode-b 
*                 |  |  |  |  |  |  |  |  |  |  |  common-anode
*                 |  |  |  |  |  |  |  |  |  |  |  |       
.SUBCKT HDSP_8600 2  3  4  5  6  7  11 12 13 14 15 17

DA1   4  2 dHDSP_8600
DB1   4 15 dHDSP_8600
DC1   4 13 dHDSP_8600
DD1   4 11 dHDSP_8600
DE1   4  5 dHDSP_8600
DF1   4  3 dHDSP_8600
DG1   4 14 dHDSP_8600
DDP1  4  7 dHDSP_8600

DA2   6  2 dHDSP_8600
DB2   6 15 dHDSP_8600
DC2   6 13 dHDSP_8600
DD2   6 11 dHDSP_8600
DE2   6  5 dHDSP_8600
DF2   6  3 dHDSP_8600
DG2   6 14 dHDSP_8600
DDP2  6  7 dHDSP_8600

DA3  12  2 dHDSP_8600
DB3  12 15 dHDSP_8600
DC3  12 13 dHDSP_8600
DD3  12 11 dHDSP_8600
DE3  12  5 dHDSP_8600
DF3  12  3 dHDSP_8600
DG3  12 14 dHDSP_8600
DDP3 12  7 dHDSP_8600

DA4  17  2 dHDSP_8600
DB4  17 15 dHDSP_8600
DC4  17 13 dHDSP_8600
DD4  17 11 dHDSP_8600
DE4  17  5 dHDSP_8600
DF4  17  3 dHDSP_8600
DG4  17 14 dHDSP_8600
DDP4 17  7 dHDSP_8600

.MODEL dHDSP_8600 D
+ (  
+     IS = 3.97670539E-22 
+      N = 1.67603447 
+     RS = 9.10910000 
+     BV = 50
+    IBV = 100u 
+ )   

.ENDS HDSP_8600
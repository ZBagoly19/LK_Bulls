*  
* Diode Model Produced by Altium Ltd  
* Date:  7-Apr-2004 
*  
* Manufacturer: Agilent  
* Component Name: HDSP-H101  
*  
* Parameters derived from information available in data sheet.  
* 
*                 cathode-e
*                 |  cathode-d
*                 |  |  common-anode
*                 |  |  |  cathode-c
*                 |  |  |  |  cathode-DP
*                 |  |  |  |  |  cathode-b
*                 |  |  |  |  |  |  cathode-a
*                 |  |  |  |  |  |  |  common-anode
*                 |  |  |  |  |  |  |  |  cathode-f
*                 |  |  |  |  |  |  |  |  |  cathode-g
*                 |  |  |  |  |  |  |  |  |  |  
.SUBCKT HDSP_H101 1  2  3  4  5  6  7  8  9  10

DA1  3  7  dHDSP_H101
DB1  3  6  dHDSP_H101
DC1  3  4  dHDSP_H101
DD1  3  2  dHDSP_H101
DE1  3  1  dHDSP_H101
DF1  3  9  dHDSP_H101
DG1  3 10  dHDSP_H101
DDP1 3  5  dHDSP_H101

DA2  8  7  dHDSP_H101
DB2  8  6  dHDSP_H101
DC2  8  4  dHDSP_H101
DD2  8  2  dHDSP_H101
DE2  8  1  dHDSP_H101
DF2  8  9  dHDSP_H101
DG2  8 10  dHDSP_H101
DDP2 8  5  dHDSP_H101

.MODEL dHDSP_H101 D
+ (  
+    IS  = 2.08276754E-16 
+     N  = 2.17799178 
+    RS  = 0.50892350
+    BV  = 14.25
+   IBV  = 100u
+ )  

.ENDS HDSP_H101
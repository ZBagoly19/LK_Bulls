*  
* Diode Model Produced by Altium Ltd  
* Date:  10-Mar-2004 
*  
* Manufacturer: Agilent  
* Component Name: HDSP-303Y  
*  
* Parameters derived from information available in data sheet.  
*
*                 anode-G
*                 |  anode-F
*                 |  |  comon-cathode
*                 |  |  |  anode-E
*                 |  |  |  |  anode-D
*                 |  |  |  |  |  anode-DP
*                 |  |  |  |  |  |  anode-C
*                 |  |  |  |  |  |  |  comon-cathode
*                 |  |  |  |  |  |  |  |  anode-B
*                 |  |  |  |  |  |  |  |  |  anode-A
*                 |  |  |  |  |  |  |  |  |  |  
.SUBCKT HDSP_303Y 1  2  3  4  5  6  7  8  9  10

DA1  10  3  dHDSP_303Y
DB1   9  3  dHDSP_303Y
DC1   7  3  dHDSP_303Y
DD1   5  3  dHDSP_303Y
DE1   4  3  dHDSP_303Y
DF1   2  3  dHDSP_303Y
DG1   1  3  dHDSP_303Y
DDP1  6  3  dHDSP_303Y

DA2  10  8  dHDSP_303Y
DB2   9  8  dHDSP_303Y
DC2   7  8  dHDSP_303Y
DD2   5  8  dHDSP_303Y
DE2   4  8  dHDSP_303Y
DF2   2  8  dHDSP_303Y
DG2   1  8  dHDSP_303Y
DDP2  6  8  dHDSP_303Y

.MODEL dHDSP_303Y D
+ (  
+     IS = 3.50837838E-27 
+      N = 1.31533553 
+     RS = 7.74814597 
+     BV = 4.8 
+    IBV = 100u 
+ )  

.ENDS HDSP_303Y
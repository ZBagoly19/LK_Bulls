*  
* Diode Model Produced by Altium Ltd  
* Date:  10-Mar-2004 
*  
* Manufacturer: Agilent  
* Component Name: HDSP-F201  
*  
* Parameters derived from information available in data sheet.  
*  
*                 common-anode 
*                 |  cathode-f 
*                 |  |  cathode-g 
*                 |  |  |  cathode-e 
*                 |  |  |  |  cathode-d 
*                 |  |  |  |  |  common-anode 
*                 |  |  |  |  |  |  cathode-DP 
*                 |  |  |  |  |  |  |  cathode-c 
*                 |  |  |  |  |  |  |  |  cathode-b 
*                 |  |  |  |  |  |  |  |  |  cathode-a
*                 |  |  |  |  |  |  |  |  |  |
.SUBCKT HDSP_F201 1  2  3  4  5  6  7  8  9  10

DA1  1 10 dHDSP_F201
DB1  1  9 dHDSP_F201
DC1  1  8 dHDSP_F201
DD1  1  5 dHDSP_F201
DE1  1  4 dHDSP_F201
DF1  1  2 dHDSP_F201
DG1  1  3 dHDSP_F201
DDP1 1  7 dHDSP_F201

DA2  6 10 dHDSP_F201
DB2  6  9 dHDSP_F201
DC2  6  8 dHDSP_F201
DD2  6  5 dHDSP_F201
DE2  6  4 dHDSP_F201
DF2  6  2 dHDSP_F201
DG2  6  3 dHDSP_F201
DDP2 6  7 dHDSP_F201

.MODEL dHDSP_F201 D
+ (  
+     IS = 3.04174763E-24 
+      N = 1.23122391 
+     RS = 24.19303791 
+     BV = 30
+    IBV = 100u 
+ )  

.ENDS HDSP_F201
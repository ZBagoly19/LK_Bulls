*  
* Diode Model Produced by Altium Ltd  
* Date:  3-May-2004 
*  
* Manufacturer: Renesas  
* Component Name: HDSP-7801  
*  
* Parameters derived from information available in data sheet.  
* 
*                 common-anode
*                 |  cathode-f
*                 |  |  cathode-g
*                 |  |  |  cathode-e
*                 |  |  |  |  cathode-d
*                 |  |  |  |  |  common-anode
*                 |  |  |  |  |  |  cathode-DP
*                 |  |  |  |  |  |  |  cathode-c
*                 |  |  |  |  |  |  |  |  cathode-b
*                 |  |  |  |  |  |  |  |  |  cathode-a
*                 |  |  |  |  |  |  |  |  |  |
.SUBCKT HDSP_7801 1  2  3  4  5  6  7  8  9  10

DA1  1  10  dHDSP_7801
DB1  1   9  dHDSP_7801
DC1  1   8  dHDSP_7801
DD1  1   5  dHDSP_7801
DE1  1   4  dHDSP_7801
DF1  1   2  dHDSP_7801
DG1  1   3  dHDSP_7801
DDP1 1   7  dHDSP_7801

DA2  6  10  dHDSP_7801
DB2  6   9  dHDSP_7801
DC2  6   8  dHDSP_7801
DD2  6   5  dHDSP_7801
DE2  6   4  dHDSP_7801
DF2  6   2  dHDSP_7801
DG2  6   3  dHDSP_7801
DDP2 6   7  dHDSP_7801

.MODEL dHDSP_7801 D
+ (  
+     IS = 1.61114016E-27 
+      N = 1.30291189 
+     RS = 12.83456794 
+     BV = 50 
+    IBV = 100u 
+ )  

.ENDS HDSP_7801
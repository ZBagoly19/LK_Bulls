*  
* Diode Model Produced by Altium Ltd  
* Date:  10-Mar-2004 
*  
* Manufacturer: Agilent  
* Component Name: HDSP-U301  
*  
* Parameters derived from information available in data sheet.  
*  
*                  cathode-a 
*                  |  cathode-f 
*                  |  |  cathode-g 
*                  |  |  |  cathode-e 
*                  |  |  |  |  cathode-d 
*                  |  |  |  |  |  cathode-DP 
*                  |  |  |  |  |  |  anode-DP 
*                  |  |  |  |  |  |  |  cathode-c 
*                  |  |  |  |  |  |  |  |  common-anode 
*                  |  |  |  |  |  |  |  |  |  cathode-b
*                  |  |  |  |  |  |  |  |  |  |
.SUBCKT HDSP_U301 1  2  3  4  5  6  7  8  9  10

D1  9  1 dHDSP_U301
D2  9  2 dHDSP_U301
D3  9  3 dHDSP_U301
D4  9  4 dHDSP_U301
D5  9  5 dHDSP_U301
D6  7  6 dHDSP_U301
D7  9  8 dHDSP_U301
D8  9 10 dHDSP_U301

.MODEL dHDSP_U301 D
+ (  
+     IS = 6.04055825E-18 
+      N = 1.90788337 
+     RS = 23.52447762 
+     BV = 40
+    IBV = 100u 
+ )  

.ENDS HDSP_U301
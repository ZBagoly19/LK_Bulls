*  
* Diode Model Produced by Altium Ltd  
* Date:  7-Apr-2004 
*  
* Manufacturer: Agilent  
* Component Name: HDSP-316L  
*  
* Parameters derived from information available in data sheet.  
* 
*                 g - anode
*                 |  f - anode
*                 |  |  common-cathode
*                 |  |  |  e - anode
*                 |  |  |  |  d - anode
*                 |  |  |  |  |  DP - anode
*                 |  |  |  |  |  |  c - anode
*                 |  |  |  |  |  |  |  common-cathode
*                 |  |  |  |  |  |  |  |  b - anode
*                 |  |  |  |  |  |  |  |  |  a - anode
*                 |  |  |  |  |  |  |  |  |  | 
.SUBCKT HDSP_316L 1  2  3  4  5  6  7  8  9  10

DA1  10 3 dHDSP_316L
DB1   9 3 dHDSP_316L
DC1   7 3 dHDSP_316L
DD1   5 3 dHDSP_316L
DE1   4 3 dHDSP_316L
DF1   2 3 dHDSP_316L
DG1   1 3 dHDSP_316L
DDP1  6 3 dHDSP_316L

DA2  10 8 dHDSP_316L
DB2   9 8 dHDSP_316L
DC2   7 8 dHDSP_316L
DD2   5 8 dHDSP_316L
DE2   4 8 dHDSP_316L
DF2   2 8 dHDSP_316L
DG2   1 8 dHDSP_316L
DDP2  6 8 dHDSP_316L

.MODEL dHDSP_316L D
+ (  
+     IS = 1.84086967E-50 
+      N = 0.55445364 
+     RS = 251.75
+     BV = 30
+    IBV = 100u 
+ )  

.ENDS HDSP_316L
*  
* Diode Model Produced by Altium Ltd  
* Date:  6-Apr-2004 
*  
* Manufacturer: Agilent  
* Component Name: HDSP-5603  
*  
* Parameters derived from information available in data sheet.  
* 
*                 anode-e
*                 |  anode-d
*                 |  |  common-cathode
*                 |  |  |  anode-c
*                 |  |  |  |  anode-DP
*                 |  |  |  |  |  anode-b
*                 |  |  |  |  |  |  anode-a
*                 |  |  |  |  |  |  |  common-cathode
*                 |  |  |  |  |  |  |  |  anode-f
*                 |  |  |  |  |  |  |  |  |  anode-g
*                 |  |  |  |  |  |  |  |  |  | 
.SUBCKT HDSP_5603 1  2  3  4  5  6  7  8  9  10

DA1   7 3 dHDSP_5603
DB1   6 3 dHDSP_5603
DC1   4 3 dHDSP_5603
DD1   2 3 dHDSP_5603
DE1   1 3 dHDSP_5603
DF1   9 3 dHDSP_5603
DG1  10 3 dHDSP_5603
DDP1  5 3 dHDSP_5603

DA2   7 8 dHDSP_5603
DB2   6 8 dHDSP_5603
DC2   4 8 dHDSP_5603
DD2   2 8 dHDSP_5603
DE2   1 8 dHDSP_5603
DF2   9 8 dHDSP_5603
DG2  10 8 dHDSP_5603
DDP2  5 8 dHDSP_5603

.MODEL dHDSP_5603 D
+ (  
+     IS = 1.61114016E-27 
+      N = 1.30291189 
+     RS = 12.83456794 
+     BV = 50 
+    IBV = 100u 
+ )

.ENDS HDSP_5603
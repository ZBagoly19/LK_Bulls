*  
* Diode Model Produced by Altium Ltd  
* Date:  3-May-2004 
*  
* Manufacturer: Renesas  
* Component Name: HDSP-7404  
*  
* Parameters derived from information available in data sheet.  
* 
*                 anode-colon
*                 |  anode-f
*                 |  |  anode-g
*                 |  |  |  anode-e
*                 |  |  |  |  anode-d
*                 |  |  |  |  |  common-cathode
*                 |  |  |  |  |  |  anode-DP
*                 |  |  |  |  |  |  |  anode-c
*                 |  |  |  |  |  |  |  |  anode-b
*                 |  |  |  |  |  |  |  |  |  anode-a
*                 |  |  |  |  |  |  |  |  |  |
.SUBCKT HDSP_7404 1  2  3  4  5  6  7  8  9  10

DA  10  6  dHDSP_7404
DB   9  6  dHDSP_7404
DC   8  6  dHDSP_7404
DD   5  6  dHDSP_7404
DE   4  6  dHDSP_7404
DF   2  6  dHDSP_7404
DG   3  6  dHDSP_7404
DDP  7  6  dHDSP_7404
DCL  1  6  dHDSP_7404

.MODEL dHDSP_7404 D
+ (  
+    IS = 2.77296438E-23 
+    N  = 1.39205436 
+    RS = 25.13253104 
+    BV = 45.00000000 
+    IBV = 100u 
+ )  

.ENDS HDSP_7404
*  
* Diode Model Produced by Altium Ltd  
* Date:  10-Mar-2004 
*  
* Manufacturer: Agilent  
* Component Name: HDSP-301G  
*  
* Parameters derived from information available in data sheet.  
*
*                 cathode-G
*                 |  cathode-F
*                 |  |  comon-anode
*                 |  |  |  cathode-E
*                 |  |  |  |  cathode-D
*                 |  |  |  |  |  cathode-DP
*                 |  |  |  |  |  |  cathode-C
*                 |  |  |  |  |  |  |  comon-anode
*                 |  |  |  |  |  |  |  |  cathode-B
*                 |  |  |  |  |  |  |  |  |  cathode-A
*                 |  |  |  |  |  |  |  |  |  |  
.SUBCKT HDSP_301G 1  2  3  4  5  6  7  8  9  10

DA1  3  10 dHDSP_301G
DB1  3   9 dHDSP_301G
DC1  3   7 dHDSP_301G
DD1  3   5 dHDSP_301G
DE1  3   4 dHDSP_301G
DF1  3   2 dHDSP_301G
DG1  3   1 dHDSP_301G
DDP1 3   6 dHDSP_301G

DA2  8  10 dHDSP_301G
DB2  8   9 dHDSP_301G
DC2  8   7 dHDSP_301G
DD2  8   5 dHDSP_301G
DE2  8   4 dHDSP_301G
DF2  8   2 dHDSP_301G
DG2  8   1 dHDSP_301G
DDP2 8   6 dHDSP_301G

.MODEL dHDSP_301G D
+ (  
+     IS = 3.14401041E-29 
+      N = 1.25233679 
+     RS = 9.99993505 
+     BV = 4.8 
+    IBV = 100u 
+ )  

.ENDS HDSP_301G
*  
* Diode Model Produced by Altium Ltd  
* Date:  10-Mar-2004 
*  
* Manufacturer: Agilent  
* Component Name: HDSP-331E  
*  
* Parameters derived from information available in data sheet.  
*  
*                 cathode-A
*                 |  cathode-F
*                 |  |  common anode
*                 |  |  |  cathode-L.DP
*                 |  |  |  |  cathode-E
*                 |  |  |  |  |  cathode-D
*                 |  |  |  |  |  |  cathode-R.DP
*                 |  |  |  |  |  |  |  cathode-C
*                 |  |  |  |  |  |  |  |  cathode-G
*                 |  |  |  |  |  |  |  |  |  cathode-B
*                 |  |  |  |  |  |  |  |  |  |  common anode
*                 |  |  |  |  |  |  |  |  |  |  |
.SUBCKT HDSP_331E 1  2  3  6  7  8  9  10 11 13 14

DA1  3  1 dHDSP_331E
DB1  3 13 dHDSP_331E
DC1  3 10 dHDSP_331E
DD1  3  8 dHDSP_331E
DE1  3  7 dHDSP_331E
DF1  3  2 dHDSP_331E
DG1  3 11 dHDSP_331E
DL1  3  6 dHDSP_331E
DR1  3  9 dHDSP_331E

DA2 14  1 dHDSP_331E
DB2 14 13 dHDSP_331E
DC2 14 10 dHDSP_331E
DD2 14  8 dHDSP_331E
DE2 14  7 dHDSP_331E
DF2 14  2 dHDSP_331E
DG2 14 11 dHDSP_331E
DL2 14  6 dHDSP_331E
DR2 14  9 dHDSP_331E

.MODEL dHDSP_331E D
+ (  
+     IS = 1.09624963E-17 
+      N = 2.02670503 
+     RS = 12.20248005 
+     BV = 4.8
+    IBV = 100u 
+ )  

.ENDS HDSP_331E
*  
* Diode Model Produced by Altium Ltd  
* Date:  10-Mar-2004 
*  
* Manufacturer: Agilent  
* Component Name: HDSP-511E  
*  
* Parameters derived from information available in data sheet.  
*  
*                 cathode-e 
*                 |  cathode-d 
*                 |  |  common-anode 
*                 |  |  |  cathode-c 
*                 |  |  |  |  cathode-DP 
*                 |  |  |  |  |  cathode-b 
*                 |  |  |  |  |  |  cathode-a 
*                 |  |  |  |  |  |  |  common-anode 
*                 |  |  |  |  |  |  |  |  cathode-f 
*                 |  |  |  |  |  |  |  |  |  cathode-g
*                 |  |  |  |  |  |  |  |  |  |
.SUBCKT HDSP_511E 1  2  3  4  5  6  7  8  9  10

DA1 3  7 dHDSP_511E
DB1 3  6 dHDSP_511E
DC1 3  4 dHDSP_511E
DD1 3  2 dHDSP_511E
DE1 3  1 dHDSP_511E
DF1 3  9 dHDSP_511E
DG1 3 10 dHDSP_511E

DA2 8  7 dHDSP_511E
DB2 8  6 dHDSP_511E
DC2 8  4 dHDSP_511E
DD2 8  2 dHDSP_511E
DE2 8  1 dHDSP_511E
DF2 8  9 dHDSP_511E
DG2 8 10 dHDSP_511E

.MODEL dHDSP_511E D
+ (  
+     IS = 6.44208414E-14 
+      N = 2.73863792 
+     RS = 11.58628790 
+     BV = 4.5
+    IBV = 100u 
+ )  

.ENDS HDSP_511E
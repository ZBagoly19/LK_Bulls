*  
* Diode Model Produced by Altium Ltd  
* Date:  6-Apr-2004 
*  
* Manufacturer: Agilent  
* Component Name: HDSP-5703  
*  
* Parameters derived from information available in data sheet.  
* 
*                 anode-e
*                 |  anode-d
*                 |  |  common-cathode
*                 |  |  |  anode-c
*                 |  |  |  |  anode-DP
*                 |  |  |  |  |  anode-b
*                 |  |  |  |  |  |  anode-a
*                 |  |  |  |  |  |  |  common-cathode
*                 |  |  |  |  |  |  |  |  anode-f
*                 |  |  |  |  |  |  |  |  |  anode-g
*                 |  |  |  |  |  |  |  |  |  | 
.SUBCKT HDSP_5703 1  2  3  4  5  6  7  8  9  10

DA1   7 3 dHDSP_5703
DB1   6 3 dHDSP_5703
DC1   4 3 dHDSP_5703
DD1   2 3 dHDSP_5703
DE1   1 3 dHDSP_5703
DF1   9 3 dHDSP_5703
DG1  10 3 dHDSP_5703
DDP1  5 3 dHDSP_5703

DA2   7 8 dHDSP_5703
DB2   6 8 dHDSP_5703
DC2   4 8 dHDSP_5703
DD2   2 8 dHDSP_5703
DE2   1 8 dHDSP_5703
DF2   9 8 dHDSP_5703
DG2  10 8 dHDSP_5703
DDP2  5 8 dHDSP_5703

.MODEL dHDSP_5703 D
+ (  
+     IS = 1.82902372E-24 
+      N = 1.34581490 
+     RS = 23.36447097 
+     BV = 40 
+    IBV = 100u 
+ )  

.ENDS HDSP_5703
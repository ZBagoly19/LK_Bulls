*  
* Diode Model Produced by Altium Ltd  
* Date:  10-Mar-2004 
*  
* Manufacturer: Agilent  
* Component Name: HDSP-F401  
*  
* Parameters derived from information available in data sheet.  
*  
*                 common-anode 
*                 |  cathode-f 
*                 |  |  cathode-g 
*                 |  |  |  cathode-e 
*                 |  |  |  |  cathode-d 
*                 |  |  |  |  |  common-anode 
*                 |  |  |  |  |  |  cathode-DP 
*                 |  |  |  |  |  |  |  cathode-c 
*                 |  |  |  |  |  |  |  |  cathode-b 
*                 |  |  |  |  |  |  |  |  |  cathode-a
*                 |  |  |  |  |  |  |  |  |  |
.SUBCKT HDSP_F401 1  2  3  4  5  6  7  8  9  10

DA1  1 10 dHDSP_F401
DB1  1  9 dHDSP_F401
DC1  1  8 dHDSP_F401
DD1  1  5 dHDSP_F401
DE1  1  4 dHDSP_F401
DF1  1  2 dHDSP_F401
DG1  1  3 dHDSP_F401
DDP1 1  7 dHDSP_F401

DA2  6 10 dHDSP_F401
DB2  6  9 dHDSP_F401
DC2  6  8 dHDSP_F401
DD2  6  5 dHDSP_F401
DE2  6  4 dHDSP_F401
DF2  6  2 dHDSP_F401
DG2  6  3 dHDSP_F401
DDP2 6  7 dHDSP_F401

.MODEL dHDSP_F401 D
+ (  
+     IS = 3.04174763E-24 
+      N = 1.23122391 
+     RS = 24.19303791 
+     BV = 30
+    IBV = 100u 
+ )  

.ENDS HDSP_F401
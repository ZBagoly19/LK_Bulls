*  
* Diode Model Produced by Altium Ltd  
* Date:  7-Apr-2004 
*  
* Manufacturer: Agilent  
* Component Name: HDSP-A901  
*  
* Parameters derived from information available in data sheet.  
*  
*                 common-anode
*                 |  cathode-f
*                 |  |  cathode-g
*                 |  |  |  cathode-e
*                 |  |  |  |  cathode-d
*                 |  |  |  |  |  common-anode
*                 |  |  |  |  |  |  cathode-DP
*                 |  |  |  |  |  |  |  cathode-c
*                 |  |  |  |  |  |  |  |  cathode-b
*                 |  |  |  |  |  |  |  |  |  cathode-a
*                 |  |  |  |  |  |  |  |  |  |
.SUBCKT HDSP_A901 1  2  3  4  5  6  7  8  9  10

DA1  1  10 dHDSP_A901
DB1  1   9 dHDSP_A901
DC1  1   8 dHDSP_A901
DD1  1   5 dHDSP_A901
DE1  1   4 dHDSP_A901
DF1  1   2 dHDSP_A901
DG1  1   3 dHDSP_A901
DDP1 1   7 dHDSP_A901

DA2  6  10 dHDSP_A901
DB2  6   9 dHDSP_A901
DC2  6   8 dHDSP_A901
DD2  6   5 dHDSP_A901
DE2  6   4 dHDSP_A901
DF2  6   2 dHDSP_A901
DG2  6   3 dHDSP_A901
DDP2 6   7 dHDSP_A901

.MODEL dHDSP_A901 D
+ (  
+     IS = 1.37135099E-36 
+      N = 0.94257009 
+     RS = 17.99091536 
+     BV = 30
+    IBV = 100u 
+ ) 

.ENDS HDSP_A901
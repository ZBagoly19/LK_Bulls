*  
* Diode Model Produced by Altium Ltd  
* Date:  10-Mar-2004 
*  
* Manufacturer: Agilent  
* Component Name: HDSP-511A  
*  
* Parameters derived from information available in data sheet.  
*  
*                 cathode-e 
*                 |  cathode-d 
*                 |  |  common-anode 
*                 |  |  |  cathode-c 
*                 |  |  |  |  cathode-DP 
*                 |  |  |  |  |  cathode-b 
*                 |  |  |  |  |  |  cathode-a 
*                 |  |  |  |  |  |  |  common-anode 
*                 |  |  |  |  |  |  |  |  cathode-f 
*                 |  |  |  |  |  |  |  |  |  cathode-g
*                 |  |  |  |  |  |  |  |  |  |
.SUBCKT HDSP_511A 1  2  3  4  5  6  7  8  9  10

DA1 3  7 dHDSP_511A
DB1 3  6 dHDSP_511A
DC1 3  4 dHDSP_511A
DD1 3  2 dHDSP_511A
DE1 3  1 dHDSP_511A
DF1 3  9 dHDSP_511A
DG1 3 10 dHDSP_511A

DA2 8  7 dHDSP_511A
DB2 8  6 dHDSP_511A
DC2 8  4 dHDSP_511A
DD2 8  2 dHDSP_511A
DE2 8  1 dHDSP_511A
DF2 8  9 dHDSP_511A
DG2 8 10 dHDSP_511A

.MODEL dHDSP_511A D
+ (  
+    IS  = 4.92088043E-22 
+     N  = 1.51994259 
+    RS  = 3.79496255
+    BV  = 4.5
+   IBV  = 100u 
+ )  

.ENDS HDSP_511A
*  
* Diode Model Produced by Altium Ltd  
* Date:  10-Mar-2004 
*  
* Manufacturer: Agilent  
* Component Name: HDSP-311G  
*  
* Parameters derived from information available in data sheet.  
* 
*                 cathode-A 
*                 |  cathode-F 
*                 |  |  common-anode 
*                 |  |  |  cathode-E 
*                 |  |  |  |  cathode-D 
*                 |  |  |  |  |  cathode-DP 
*                 |  |  |  |  |  |  cathode-C 
*                 |  |  |  |  |  |  |  cathode-G 
*                 |  |  |  |  |  |  |  |  cathode-B 
*                 |  |  |  |  |  |  |  |  |  common-anode
*                 |  |  |  |  |  |  |  |  |  |
.SUBCKT HDSP_311G 1  2  3  7  8  9  10 11 13 14

DA1   3  1 dHDSP_311G
DB1   3 13 dHDSP_311G
DC1   3 10 dHDSP_311G
DD1   3  8 dHDSP_311G
DE1   3  7 dHDSP_311G
DF1   3  2 dHDSP_311G
DG1   3 11 dHDSP_311G
DDP1  3  9 dHDSP_311G

DA2  14  1 dHDSP_311G
DB2  14 13 dHDSP_311G
DC2  14 10 dHDSP_311G
DD2  14  8 dHDSP_311G
DE2  14  7 dHDSP_311G
DF2  14  2 dHDSP_311G
DG2  14 11 dHDSP_311G
DDP2 14  9 dHDSP_311G

.MODEL dHDSP_311G D
+ (  
+     IS = 1.61114016E-27 
+      N = 1.30291189 
+     RS = 12.83456794 
+     BV = 50 
+    IBV = 100u 
+ )  

.ENDS HDSP_311G
*  
* Diode Model Produced by Altium Ltd  
* Date:  7-Apr-2004 
*  
* Manufacturer: Agilent  
* Component Name: HDSP-4603  
*  
* Parameters derived from information available in data sheet.  
* 
*                 anode-a
*                 |  anode-f
*                 |  |  common-cathode
*                 |  |  |  anode-e
*                 |  |  |  |  anode-d
*                 |  |  |  |  |  anode-DP
*                 |  |  |  |  |  |  anode-c
*                 |  |  |  |  |  |  |  anode-g
*                 |  |  |  |  |  |  |  |  anode-b
*                 |  |  |  |  |  |  |  |  |  common-cathode
*                 |  |  |  |  |  |  |  |  |  |
.SUBCKT HDSP_4603 1  2  3  7  8  9  10 11 13 14

DA1   1  3 dHDSP_4603
DB1  13  3 dHDSP_4603
DC1  10  3 dHDSP_4603
DD1   8  3 dHDSP_4603
DE1   7  3 dHDSP_4603
DF1   2  3 dHDSP_4603
DG1  11  3 dHDSP_4603
DDP1  9  3 dHDSP_4603

DA2   1 14 dHDSP_4603
DB2  13 14 dHDSP_4603
DC2  10 14 dHDSP_4603
DD2   8 14 dHDSP_4603
DE2   7 14 dHDSP_4603
DF2   2 14 dHDSP_4603
DG2  11 14 dHDSP_4603
DDP2  9 14 dHDSP_4603

.MODEL dHDSP_4603 D
+ (  
+     IS = 1.61114016E-27 
+      N = 1.30291189 
+     RS = 12.83456794 
+     BV = 50 
+    IBV = 100u 
+ )  

.ENDS HDSP_4603
*  
* Diode Model Produced by Altium Ltd  
* Date:  10-Mar-2004 
*  
* Manufacturer: Agilent  
* Component Name: HDSP-F151  
*  
* Parameters derived from information available in data sheet.  
*  
*                 common-anode 
*                 |  cathode-f 
*                 |  |  cathode-g 
*                 |  |  |  cathode-e 
*                 |  |  |  |  cathode-d 
*                 |  |  |  |  |  common-anode 
*                 |  |  |  |  |  |  cathode-DP 
*                 |  |  |  |  |  |  |  cathode-c 
*                 |  |  |  |  |  |  |  |  cathode-b 
*                 |  |  |  |  |  |  |  |  |  cathode-a
*                 |  |  |  |  |  |  |  |  |  |
.SUBCKT HDSP_F151 1  2  3  4  5  6  7  8  9  10

DA1  1 10 dHDSP_F151
DB1  1  9 dHDSP_F151
DC1  1  8 dHDSP_F151
DD1  1  5 dHDSP_F151
DE1  1  4 dHDSP_F151
DF1  1  2 dHDSP_F151
DG1  1  3 dHDSP_F151
DDP1 1  7 dHDSP_F151

DA2  6 10 dHDSP_F151
DB2  6  9 dHDSP_F151
DC2  6  8 dHDSP_F151
DD2  6  5 dHDSP_F151
DE2  6  4 dHDSP_F151
DF2  6  2 dHDSP_F151
DG2  6  3 dHDSP_F151
DDP2 6  7 dHDSP_F151

.MODEL dHDSP_F151 D
+ (  
+    IS  = 1.31055154E-15 
+     N  = 2.20660855 
+    RS  = 1.60736539 
+    BV  = 14.25
+   IBV  = 100u
+ )  

.ENDS HDSP_F151
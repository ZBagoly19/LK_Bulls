*  
* Diode Model Produced by Altium Ltd  
* Date:  7-Apr-2004 
*  
* Manufacturer: Agilent  
* Component Name: HDSP-E103  
*  
* Parameters derived from information available in data sheet.  
*  
*                 anode-a
*                 |  anode-f
*                 |  |  common-cathode
*                 |  |  |  anode-e
*                 |  |  |  |  anode-d
*                 |  |  |  |  |  anode-DP
*                 |  |  |  |  |  |  anode-c
*                 |  |  |  |  |  |  |  anode-g
*                 |  |  |  |  |  |  |  |  anode-b
*                 |  |  |  |  |  |  |  |  |  common-cathode
*                 |  |  |  |  |  |  |  |  |  |
.SUBCKT HDSP_E103 1  2  3  7  8  9  10 11 13 14

DA1   1   3 dHDSP_E103
DB1  13   3 dHDSP_E103
DC1  10   3 dHDSP_E103
DD1   8   3 dHDSP_E103
DE1   7   3 dHDSP_E103
DF1   2   3 dHDSP_E103
DG1  11   3 dHDSP_E103
DDP1  9   3 dHDSP_E103

DA2   1  14 dHDSP_E103
DB2  13  14 dHDSP_E103
DC2  10  14 dHDSP_E103
DD2   8  14 dHDSP_E103
DE2   7  14 dHDSP_E103
DF2   2  14 dHDSP_E103
DG2  11  14 dHDSP_E103
DDP2  9  14 dHDSP_E103

.MODEL dHDSP_E103 D
+ (  
+    IS  = 2.08276754E-16 
+     N  = 2.17799178 
+    RS  = 0.50892350
+    BV  = 14.25
+   IBV  = 100u
+ )

.ENDS HDSP_E103
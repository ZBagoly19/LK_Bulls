*  
* Diode Model Produced by Altium Ltd  
* Date:  7-Apr-2004 
*  
* Manufacturer: Agilent  
* Component Name: HDSP-316G  
*  
* Parameters derived from information available in data sheet.  
* 
*                 g - anode
*                 |  f - anode
*                 |  |  common-cathode
*                 |  |  |  e - anode
*                 |  |  |  |  d - anode
*                 |  |  |  |  |  DP - anode
*                 |  |  |  |  |  |  c - anode
*                 |  |  |  |  |  |  |  common-cathode
*                 |  |  |  |  |  |  |  |  b - anode
*                 |  |  |  |  |  |  |  |  |  a - anode
*                 |  |  |  |  |  |  |  |  |  | 
.SUBCKT HDSP_316G 1  2  3  4  5  6  7  8  9  10

DA1  10 3 dHDSP_316G
DB1   9 3 dHDSP_316G
DC1   7 3 dHDSP_316G
DD1   5 3 dHDSP_316G
DE1   4 3 dHDSP_316G
DF1   2 3 dHDSP_316G
DG1   1 3 dHDSP_316G
DDP1  6 3 dHDSP_316G

DA2  10 8 dHDSP_316G
DB2   9 8 dHDSP_316G
DC2   7 8 dHDSP_316G
DD2   5 8 dHDSP_316G
DE2   4 8 dHDSP_316G
DF2   2 8 dHDSP_316G
DG2   1 8 dHDSP_316G
DDP2  6 8 dHDSP_316G

.MODEL dHDSP_316G D
+ (  
+     IS = 1.61114016E-27 
+      N = 1.30291189 
+     RS = 12.83456794 
+     BV = 50 
+    IBV = 100u 
+ )  

.ENDS HDSP_316G
*  
* Diode Model Produced by Altium Ltd  
* Date:  10-Mar-2004 
*  
* Manufacturer: Agilent  
* Component Name: HDSP-H111  
*  
* Parameters derived from information available in data sheet.  
* 
*                 cathode-e
*                 |  cathode-d
*                 |  |  common-anode
*                 |  |  |  cathode-c
*                 |  |  |  |  cathode-DP
*                 |  |  |  |  |  cathode-b
*                 |  |  |  |  |  |  cathode-a
*                 |  |  |  |  |  |  |  common-anode
*                 |  |  |  |  |  |  |  |  cathode-f
*                 |  |  |  |  |  |  |  |  |  cathode-g
*                 |  |  |  |  |  |  |  |  |  | 
.SUBCKT HDSP_H111 1  2  3  4  5  6  7  8  9  10

DA1   3  7  dHDSP_H111
DB1   3  6  dHDSP_H111
DC1   3  4  dHDSP_H111
DD1   3  2  dHDSP_H111
DE1   3  1  dHDSP_H111
DF1   3  9  dHDSP_H111
DG1   3 10  dHDSP_H111
DDP1  3  5  dHDSP_H111

DA2   8  7  dHDSP_H111
DB2   8  6  dHDSP_H111
DC2   8  4  dHDSP_H111
DD2   8  2  dHDSP_H111
DE2   8  1  dHDSP_H111
DF2   8  9  dHDSP_H111
DG2   8 10  dHDSP_H111
DDP2  8  5  dHDSP_H111

.MODEL dHDSP_H111 D
+ (  
+    IS  = 2.08276754E-16 
+     N  = 2.17799178 
+    RS  = 0.50892350
+    BV  = 14.25
+   IBV  = 100u
+ )  

.ENDS HDSP_H111
*  
* Diode Model Produced by Altium Ltd  
* Date:  7-Apr-2004 
*  
* Manufacturer: Agilent  
* Component Name: HDSP-3351  
*  
* Parameters derived from information available in data sheet.  
*  
*                 cathode-a
*                 |  cathode-f
*                 |  |  common-anode
*                 |  |  |  cathode-e
*                 |  |  |  |  cathode-d
*                 |  |  |  |  |  cathode-DP
*                 |  |  |  |  |  |  cathode-c
*                 |  |  |  |  |  |  |  cathode-g
*                 |  |  |  |  |  |  |  |  cathode-b
*                 |  |  |  |  |  |  |  |  |  common-anode
*                 |  |  |  |  |  |  |  |  |  |
.SUBCKT HDSP_3351 1  2  3  7  8  9  10 11 13 14

DA1   3   1 dHDSP_3351
DB1   3  13 dHDSP_3351
DC1   3  10 dHDSP_3351
DD1   3   8 dHDSP_3351
DE1   3   7 dHDSP_3351
DF1   3   2 dHDSP_3351
DG1   3  11 dHDSP_3351
DDP1  3   9 dHDSP_3351

DA2  14   1 dHDSP_3351
DB2  14  13 dHDSP_3351
DC2  14  10 dHDSP_3351
DD2  14   8 dHDSP_3351
DE2  14   7 dHDSP_3351
DF2  14   2 dHDSP_3351
DG2  14  11 dHDSP_3351
DDP2 14   9 dHDSP_3351

.MODEL dHDSP_3351 D
+ (  
+     IS = 7.07436607E-24 
+      N = 1.24380258 
+     RS = 22.12166762 
+     BV = 30
+    IBV = 100u 
+ )  

.ENDS HDSP_3351
*  
* Diode Model Produced by Altium Ltd  
* Date:  7-Apr-2004 
*  
* Manufacturer: Agilent  
* Component Name: HDSP-5731  
*  
* Parameters derived from information available in data sheet.  
*
*                 e 
*                 |  d 
*                 |  |  common-anode
*                 |  |  |  c 
*                 |  |  |  |  DP  
*                 |  |  |  |  |  b 
*                 |  |  |  |  |  |  a 
*                 |  |  |  |  |  |  |  common-anode   
*                 |  |  |  |  |  |  |  |  f  
*                 |  |  |  |  |  |  |  |  |  g
*                 |  |  |  |  |  |  |  |  |  |  
.SUBCKT HDSP_5731 1  2  3  4  5  6  7  8  9  10

DA1  3  7 dHDSP_5731
DB1  3  6 dHDSP_5731
DC1  3  4 dHDSP_5731
DD1  3  2 dHDSP_5731
DE1  3  1 dHDSP_5731
DF1  3  9 dHDSP_5731
DG1  3 10 dHDSP_5731
DDP1 3  5 dHDSP_5731

DA2  8  7 dHDSP_5731
DB2  8  6 dHDSP_5731
DC2  8  4 dHDSP_5731
DD2  8  2 dHDSP_5731
DE2  8  1 dHDSP_5731
DF2  8  9 dHDSP_5731
DG2  8 10 dHDSP_5731
DDP2 8  5 dHDSP_5731

.MODEL dHDSP_5731 D
+ (  
+     IS = 8.07922028E-13 
+      N = 3.08151986 
+     RS = 5.65168121 
+     BV = 2.25
+    IBV = 100u 
+ )  

.ENDS HDSP_4136
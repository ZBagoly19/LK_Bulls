*  
* Diode Model Produced by Altium Ltd  
* Date:  10-Mar-2004 
*  
* Manufacturer: Agilent  
* Component Name: HDSP-563Y  
*  
* Parameters derived from information available in data sheet.  
*
*                 anode-E
*                 |  anode-D
*                 |  |  comon-cathode
*                 |  |  |  anode-C
*                 |  |  |  |  anode-DP
*                 |  |  |  |  |  anode-B
*                 |  |  |  |  |  |  anode-A
*                 |  |  |  |  |  |  |  comon-cathode
*                 |  |  |  |  |  |  |  |  anode-F
*                 |  |  |  |  |  |  |  |  |  anode-G
*                 |  |  |  |  |  |  |  |  |  |  
.SUBCKT HDSP_563Y 1  2  3  4  5  6  7  8  9  10

DA1   7  3  dHDSP_563Y
DB1   6  3  dHDSP_563Y
DC1   4  3  dHDSP_563Y
DD1   2  3  dHDSP_563Y
DE1   1  3  dHDSP_563Y
DF1   9  3  dHDSP_563Y
DG1  10  3  dHDSP_563Y
DDP1  5  3  dHDSP_563Y

DA2   7  8  dHDSP_563Y
DB2   6  8  dHDSP_563Y
DC2   4  8  dHDSP_563Y
DD2   2  8  dHDSP_563Y
DE2   1  8  dHDSP_563Y
DF2   9  8  dHDSP_563Y
DG2  10  8  dHDSP_563Y
DDP2  5  8  dHDSP_563Y

.MODEL dHDSP_563Y D
+ (  
+     IS = 3.50837838E-27 
+      N = 1.31533553 
+     RS = 7.74814597 
+     BV = 4.8 
+    IBV = 100u 
+ )  

.ENDS HDSP_563Y
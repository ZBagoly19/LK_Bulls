*  
* Diode Model Produced by Altium Ltd  
* Date:  7-Apr-2004 
*  
* Manufacturer: Agilent  
* Component Name: HDSP-N153  
*  
* Parameters derived from information available in data sheet.  
*  
*                 anode-a 
*                 |  anode-f 
*                 |  |  common-cathode 
*                 |  |  |  anode-e 
*                 |  |  |  |  common-cathode 
*                 |  |  |  |  |  anode-DP 
*                 |  |  |  |  |  |  anode-d 
*                 |  |  |  |  |  |  |  common-cathode 
*                 |  |  |  |  |  |  |  |  anode-c 
*                 |  |  |  |  |  |  |  |  |  anode-g 
*                 |  |  |  |  |  |  |  |  |  |  anode-b 
*                 |  |  |  |  |  |  |  |  |  |  |  common-cathode
*                 |  |  |  |  |  |  |  |  |  |  |  |       
.SUBCKT HDSP_N153 2  3  4  5  6  10 11 12 13 14 15 17

DA1   2  4 dHDSP_N153
DB1  15  4 dHDSP_N153
DC1  13  4 dHDSP_N153
DD1  11  4 dHDSP_N153
DE1   5  4 dHDSP_N153
DF1   3  4 dHDSP_N153
DG1  14  4 dHDSP_N153
DDP1 10  4 dHDSP_N153

DA2   2  6 dHDSP_N153
DB2  15  6 dHDSP_N153
DC2  13  6 dHDSP_N153
DD2  11  6 dHDSP_N153
DE2   5  6 dHDSP_N153
DF2   3  6 dHDSP_N153
DG2  14  6 dHDSP_N153
DDP2 10  6 dHDSP_N153

DA3   2 12 dHDSP_N153
DB3  15 12 dHDSP_N153
DC3  13 12 dHDSP_N153
DD3  11 12 dHDSP_N153
DE3   5 12 dHDSP_N153
DF3   3 12 dHDSP_N153
DG3  14 12 dHDSP_N153
DDP3 10 12 dHDSP_N153

DA4   2 17 dHDSP_N153
DB4  15 17 dHDSP_N153
DC4  13 17 dHDSP_N153
DD4  11 17 dHDSP_N153
DE4   5 17 dHDSP_N153
DF4   3 17 dHDSP_N153
DG4  14 17 dHDSP_N153
DDP4 10 17 dHDSP_N153

.MODEL dHDSP_N153 D
+ (  
+    IS = 1.72301609E-14 
+     N = 2.43230682 
+    RS = 1.67295284
+    BV = 14.25
+   IBV = 100u 
+ )  

.ENDS HDSP_N153
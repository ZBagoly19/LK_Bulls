*  
* Diode Model Produced by Altium Ltd  
* Date:  6-Apr-2004 
*  
* Manufacturer: Agilent  
* Component Name: HDSP-5523  
*  
* Parameters derived from information available in data sheet.  
* 
*                 E-anode-1
*                 |  D-anode-1
*                 |  |  C-anode-1
*                 |  |  |  DP-anode-1
*                 |  |  |  |  E-anode-1
*                 |  |  |  |  |  D-anode-2
*                 |  |  |  |  |  |  G-anode-2
*                 |  |  |  |  |  |  |  C-anode-2
*                 |  |  |  |  |  |  |  |  DP-anode-2
*                 |  |  |  |  |  |  |  |  |  B-anode-2
*                 |  |  |  |  |  |  |  |  |  |  A-anode-2
*                 |  |  |  |  |  |  |  |  |  |  |  F-anode-2
*                 |  |  |  |  |  |  |  |  |  |  |  |  common-cathode-2
*                 |  |  |  |  |  |  |  |  |  |  |  |  |  common-cathode-1
*                 |  |  |  |  |  |  |  |  |  |  |  |  |  |  B-anode-1
*                 |  |  |  |  |  |  |  |  |  |  |  |  |  |  |  A-anode-1
*                 |  |  |  |  |  |  |  |  |  |  |  |  |  |  |  |  G-anode-1
*                 |  |  |  |  |  |  |  |  |  |  |  |  |  |  |  |  |  F-anode-1
*                 |  |  |  |  |  |  |  |  |  |  |  |  |  |  |  |  |  |
.SUBCKT HDSP_5523 1  2  3  4  5  6  7  8  9  10 11 12 13 14 15 16 17 18

DA1  16  14  dHDSP_5523
DB1  15  14  dHDSP_5523
DC1   3  14  dHDSP_5523
DD1   2  14  dHDSP_5523
DE1   1  14  dHDSP_5523
DF1  18  14  dHDSP_5523
DG1  17  14  dHDSP_5523
DDP1  4  14  dHDSP_5523

DA2  11  13  dHDSP_5523
DB2  10  13  dHDSP_5523
DC2   8  13  dHDSP_5523
DD2   6  13  dHDSP_5523
DE2   5  13  dHDSP_5523
DF2  12  13  dHDSP_5523
DG2   7  13  dHDSP_5523
DDP2  9  13  dHDSP_5523

.MODEL dHDSP_5523 D
+ (  
+     IS = 3.78006861E-14 
+      N = 2.44553183 
+     RS = 19.51958310 
+     BV = 30
+    IBV = 100u 
+ )  

.ENDS HDSP_5523
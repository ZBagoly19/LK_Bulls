*  
* Diode Model Produced by Altium Ltd  
* Date:  10-Mar-2004 
*  
* Manufacturer: Agilent  
* Component Name: HDSP-U501  
*  
* Parameters derived from information available in data sheet.  
*  
*                  cathode-a 
*                  |  cathode-f 
*                  |  |  cathode-g 
*                  |  |  |  cathode-e 
*                  |  |  |  |  cathode-d 
*                  |  |  |  |  |  cathode-DP 
*                  |  |  |  |  |  |  anode-DP 
*                  |  |  |  |  |  |  |  cathode-c 
*                  |  |  |  |  |  |  |  |  common-anode 
*                  |  |  |  |  |  |  |  |  |  cathode-b
*                  |  |  |  |  |  |  |  |  |  |
.SUBCKT HDSP_U501 1  2  3  4  5  6  7  8  9  10

D1  9  1 dHDSP_U501
D2  9  2 dHDSP_U501
D3  9  3 dHDSP_U501
D4  9  4 dHDSP_U501
D5  9  5 dHDSP_U501
D6  7  6 dHDSP_U501
D7  9  8 dHDSP_U501
D8  9 10 dHDSP_U501

.MODEL dHDSP_U501 D
+ (  
+     IS = 1.61114016E-27 
+      N = 1.30291189 
+     RS = 12.83456794 
+     BV = 50 
+    IBV = 100u 
+ )  

.ENDS HDSP_U501
*  
* Diode Model Produced by Altium Ltd  
* Date:  7-Apr-2004 
*  
* Manufacturer: Agilent  
* Component Name: HDSP-516E  
*  
* Parameters derived from information available in data sheet.  
* 
*                 e - anode
*                 |  d - anode
*                 |  |  common-cathode
*                 |  |  |  c - anode
*                 |  |  |  |  DP - anode
*                 |  |  |  |  |  b - anode
*                 |  |  |  |  |  |  a - anode
*                 |  |  |  |  |  |  |  common-cathode
*                 |  |  |  |  |  |  |  |  f - anode
*                 |  |  |  |  |  |  |  |  |  g - anode
*                 |  |  |  |  |  |  |  |  |  | 
.SUBCKT HDSP_516E 1  2  3  4  5  6  7  8  9  10

DA1   7 3 dHDSP_516E
DB1   6 3 dHDSP_516E
DC1   4 3 dHDSP_516E
DD1   2 3 dHDSP_516E
DE1   1 3 dHDSP_516E
DF1   9 3 dHDSP_516E
DG1  10 3 dHDSP_516E
DDP1  5 3 dHDSP_516E

DA2   7 8 dHDSP_516E
DB2   6 8 dHDSP_516E
DC2   4 8 dHDSP_516E
DD2   2 8 dHDSP_516E
DE2   1 8 dHDSP_516E
DF2   9 8 dHDSP_516E
DG2  10 8 dHDSP_516E
DDP2  5 8 dHDSP_516E

.MODEL dHDSP_516E D
+ (  
+     IS = 1.21481726E-49 
+      N = 0.55445364 
+     RS = 25.38287000 
+     BV = 30
+    IBV = 100u 
+ )  

.ENDS HDSP_516E
*  
* Diode Model Produced by Altium Ltd  
* Date:  10-Mar-2004 
*  
* Manufacturer: Agilent  
* Component Name: HDSP-U103  
*  
* Parameters derived from information available in data sheet.  
*  
*                  anode-a 
*                  |  anode-f 
*                  |  |  anode-g 
*                  |  |  |  anode-e 
*                  |  |  |  |  anode-d 
*                  |  |  |  |  |  cathode-DP 
*                  |  |  |  |  |  |  anode-DP 
*                  |  |  |  |  |  |  |  anode-c 
*                  |  |  |  |  |  |  |  |  common-cathode 
*                  |  |  |  |  |  |  |  |  |  anode-b
*                  |  |  |  |  |  |  |  |  |  |
.SUBCKT HDSP_U103 1  2  3  4  5  6  7  8  9  10

D1  1  9 dHDSP_U103
D2  2  9 dHDSP_U103
D3  3  9 dHDSP_U103
D4  4  9 dHDSP_U103
D5  5  9 dHDSP_U103
D6  7  6 dHDSP_U103
D7  8  9 dHDSP_U103
D8 10  9 dHDSP_U103

.MODEL dHDSP_U103 D
+ (  
+    IS  = 1.31055154E-15 
+     N  = 2.20660855 
+    RS  = 1.60736539 
+    BV  = 14.25
+   IBV  = 100u
+ )  

.ENDS HDSP_U103
*  
* Diode Model Produced by Altium Ltd  
* Date:  7-Apr-2004 
*  
* Manufacturer: Agilent  
* Component Name: HDSP-315Y  
*  
* Parameters derived from information available in data sheet.  
* 
*                 g - cathode
*                 |  f - cathode
*                 |  |  common-anode
*                 |  |  |  e - cathode
*                 |  |  |  |  d - cathode
*                 |  |  |  |  |  DP - cathode
*                 |  |  |  |  |  |  c - cathode
*                 |  |  |  |  |  |  |  common-anode
*                 |  |  |  |  |  |  |  |  b - cathode
*                 |  |  |  |  |  |  |  |  |  a - cathode
*                 |  |  |  |  |  |  |  |  |  | 
.SUBCKT HDSP_315Y 1  2  3  4  5  6  7  8  9  10

DA1  3 10 dHDSP_315Y
DB1  3  9 dHDSP_315Y
DC1  3  7 dHDSP_315Y
DD1  3  5 dHDSP_315Y
DE1  3  4 dHDSP_315Y
DF1  3  2 dHDSP_315Y
DG1  3  1 dHDSP_315Y
DDP1 3  6 dHDSP_315Y

DA2  8 10 dHDSP_315Y
DB2  8  9 dHDSP_315Y
DC2  8  7 dHDSP_315Y
DD2  8  5 dHDSP_315Y
DE2  8  4 dHDSP_315Y
DF2  8  2 dHDSP_315Y
DG2  8  1 dHDSP_315Y
DDP2 8  6 dHDSP_315Y

.MODEL dHDSP_315Y D
+ (  
+     IS = 3.94588412E-15 
+      N = 2.33201916 
+     RS = 23.30053910 
+     BV = 50 
+    IBV = 100u 
+ )  

.ENDS HDSP_315Y
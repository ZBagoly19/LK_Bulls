*  
* Diode Model Produced by Altium Ltd  
* Date:  7-Apr-2004 
*  
* Manufacturer: Agilent  
* Component Name: HDSP-516Y  
*  
* Parameters derived from information available in data sheet.  
* 
*                 e - anode
*                 |  d - anode
*                 |  |  common-cathode
*                 |  |  |  c - anode
*                 |  |  |  |  DP - anode
*                 |  |  |  |  |  b - anode
*                 |  |  |  |  |  |  a - anode
*                 |  |  |  |  |  |  |  common-cathode
*                 |  |  |  |  |  |  |  |  f - anode
*                 |  |  |  |  |  |  |  |  |  g - anode
*                 |  |  |  |  |  |  |  |  |  | 
.SUBCKT HDSP_516Y 1  2  3  4  5  6  7  8  9  10

DA1   7 3 dHDSP_516Y
DB1   6 3 dHDSP_516Y
DC1   4 3 dHDSP_516Y
DD1   2 3 dHDSP_516Y
DE1   1 3 dHDSP_516Y
DF1   9 3 dHDSP_516Y
DG1  10 3 dHDSP_516Y
DDP1  5 3 dHDSP_516Y

DA2   7 8 dHDSP_516Y
DB2   6 8 dHDSP_516Y
DC2   4 8 dHDSP_516Y
DD2   2 8 dHDSP_516Y
DE2   1 8 dHDSP_516Y
DF2   9 8 dHDSP_516Y
DG2  10 8 dHDSP_516Y
DDP2  5 8 dHDSP_516Y

.MODEL dHDSP_516Y D
+ (  
+     IS = 3.94588412E-15 
+      N = 2.33201916 
+     RS = 23.30053910 
+     BV = 50 
+    IBV = 100u 
+ )  

.ENDS HDSP_516Y
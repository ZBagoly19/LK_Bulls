*  
* Diode Model Produced by Altium Ltd  
* Date:  10-Mar-2004 
*  
* Manufacturer: Agilent  
* Component Name: HDSP-563E  
*  
* Parameters derived from information available in data sheet.  
*
*                 anode-E
*                 |  anode-D
*                 |  |  comon-cathode
*                 |  |  |  anode-C
*                 |  |  |  |  anode-DP
*                 |  |  |  |  |  anode-B
*                 |  |  |  |  |  |  anode-A
*                 |  |  |  |  |  |  |  comon-cathode
*                 |  |  |  |  |  |  |  |  anode-F
*                 |  |  |  |  |  |  |  |  |  anode-G
*                 |  |  |  |  |  |  |  |  |  |  
.SUBCKT HDSP_563E 1  2  3  4  5  6  7  8  9  10

DA1   7  3  dHDSP_563E
DB1   6  3  dHDSP_563E
DC1   4  3  dHDSP_563E
DD1   2  3  dHDSP_563E
DE1   1  3  dHDSP_563E
DF1   9  3  dHDSP_563E
DG1  10  3  dHDSP_563E
DDP1  5  3  dHDSP_563E

DA2   7  8  dHDSP_563E
DB2   6  8  dHDSP_563E
DC2   4  8  dHDSP_563E
DD2   2  8  dHDSP_563E
DE2   1  8  dHDSP_563E
DF2   9  8  dHDSP_563E
DG2  10  8  dHDSP_563E
DDP2  5  8  dHDSP_563E

.MODEL dHDSP_563E D
+ (  
+     IS = 1.37607512E-24 
+      N = 1.38335616 
+     RS = 6.06238569 
+     BV = 4.8 
+    IBV = 100u 
+ ) 

.ENDS HDSP_563E
*  
* Diode Model Produced by Altium Ltd  
* Date:  10-Mar-2004 
*  
* Manufacturer: Agilent  
* Component Name: HDSP-F301  
*  
* Parameters derived from information available in data sheet.  
*  
*                 common-anode 
*                 |  cathode-f 
*                 |  |  cathode-g 
*                 |  |  |  cathode-e 
*                 |  |  |  |  cathode-d 
*                 |  |  |  |  |  common-anode 
*                 |  |  |  |  |  |  cathode-DP 
*                 |  |  |  |  |  |  |  cathode-c 
*                 |  |  |  |  |  |  |  |  cathode-b 
*                 |  |  |  |  |  |  |  |  |  cathode-a
*                 |  |  |  |  |  |  |  |  |  |
.SUBCKT HDSP_F301 1  2  3  4  5  6  7  8  9  10

DA1  1 10 dHDSP_F301
DB1  1  9 dHDSP_F301
DC1  1  8 dHDSP_F301
DD1  1  5 dHDSP_F301
DE1  1  4 dHDSP_F301
DF1  1  2 dHDSP_F301
DG1  1  3 dHDSP_F301
DDP1 1  7 dHDSP_F301

DA2  6 10 dHDSP_F301
DB2  6  9 dHDSP_F301
DC2  6  8 dHDSP_F301
DD2  6  5 dHDSP_F301
DE2  6  4 dHDSP_F301
DF2  6  2 dHDSP_F301
DG2  6  3 dHDSP_F301
DDP2 6  7 dHDSP_F301

.MODEL dHDSP_F301 D
+ (  
+     IS = 6.04055825E-18 
+      N = 1.90788337 
+     RS = 23.52447762 
+     BV = 40
+    IBV = 100u 
+ )  

.ENDS HDSP_F301
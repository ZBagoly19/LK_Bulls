*  
* Diode Model Produced by Altium Ltd  
* Date:  7-Apr-2004 
*  
* Manufacturer: Agilent  
* Component Name: HDSP-A101  
*  
* Parameters derived from information available in data sheet.  
*  
*                 common-anode
*                 |  cathode-f
*                 |  |  cathode-g
*                 |  |  |  cathode-e
*                 |  |  |  |  cathode-d
*                 |  |  |  |  |  common-anode
*                 |  |  |  |  |  |  cathode-DP
*                 |  |  |  |  |  |  |  cathode-c
*                 |  |  |  |  |  |  |  |  cathode-b
*                 |  |  |  |  |  |  |  |  |  cathode-a
*                 |  |  |  |  |  |  |  |  |  |
.SUBCKT HDSP_A101 1  2  3  4  5  6  7  8  9  10

DA1  1  10 dHDSP_A101
DB1  1   9 dHDSP_A101
DC1  1   8 dHDSP_A101
DD1  1   5 dHDSP_A101
DE1  1   4 dHDSP_A101
DF1  1   2 dHDSP_A101
DG1  1   3 dHDSP_A101
DDP1 1   7 dHDSP_A101

DA2  6  10 dHDSP_A101
DB2  6   9 dHDSP_A101
DC2  6   8 dHDSP_A101
DD2  6   5 dHDSP_A101
DE2  6   4 dHDSP_A101
DF2  6   2 dHDSP_A101
DG2  6   3 dHDSP_A101
DDP2 6   7 dHDSP_A101

.MODEL dHDSP_A101 D
+ (  
+    IS  = 2.08276754E-16 
+     N  = 2.17799178 
+    RS  = 0.50892350
+    BV  = 14.25
+   IBV  = 100u
+ ) 

.ENDS HDSP_A101
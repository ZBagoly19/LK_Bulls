*  
* Diode Model Produced by Altium Ltd  
* Date:  6-Apr-2004 
*  
* Manufacturer: Agilent  
* Component Name: HDSP-H153  
*  
* Parameters derived from information available in data sheet.  
* 
*                 anode-e
*                 |  anode-d
*                 |  |  common-cathode
*                 |  |  |  anode-c
*                 |  |  |  |  anode-DP
*                 |  |  |  |  |  anode-b
*                 |  |  |  |  |  |  anode-a
*                 |  |  |  |  |  |  |  common-cathode
*                 |  |  |  |  |  |  |  |  anode-f
*                 |  |  |  |  |  |  |  |  |  anode-g
*                 |  |  |  |  |  |  |  |  |  | 
.SUBCKT HDSP_H153 1  2  3  4  5  6  7  8  9  10

DA1   7 3 dHDSP_H153
DB1   6 3 dHDSP_H153
DC1   4 3 dHDSP_H153
DD1   2 3 dHDSP_H153
DE1   1 3 dHDSP_H153
DF1   9 3 dHDSP_H153
DG1  10 3 dHDSP_H153
DDP1  5 3 dHDSP_H153

DA2   7 8 dHDSP_H153
DB2   6 8 dHDSP_H153
DC2   4 8 dHDSP_H153
DD2   2 8 dHDSP_H153
DE2   1 8 dHDSP_H153
DF2   9 8 dHDSP_H153
DG2  10 8 dHDSP_H153
DDP2  5 8 dHDSP_H153

.MODEL dHDSP_H153 D
+ (  
+    IS = 3.25509599E-15 
+     N = 2.27697656 
+    RS = 1.58416732
+    BV = 14.25
+   IBV = 100u
+ ) 

.ENDS HDSP_H153
*  
* Diode Model Produced by Altium Ltd  
* Date:  7-Apr-2004 
*  
* Manufacturer: Agilent  
* Component Name: HDSP-8601  
*  
* Parameters derived from information available in data sheet.  
*  
*                 cathode-a 
*                 |  cathode-f 
*                 |  |  common-anode 
*                 |  |  |  cathode-e 
*                 |  |  |  |  common-anode 
*                 |  |  |  |  |  cathode-DP 
*                 |  |  |  |  |  |  cathode-d 
*                 |  |  |  |  |  |  |  common-anode 
*                 |  |  |  |  |  |  |  |  cathode-c 
*                 |  |  |  |  |  |  |  |  |  cathode-g 
*                 |  |  |  |  |  |  |  |  |  |  cathode-b 
*                 |  |  |  |  |  |  |  |  |  |  |  common-anode
*                 |  |  |  |  |  |  |  |  |  |  |  |       
.SUBCKT HDSP_8601 2  3  4  5  6  10 11 12 13 14 15 17

DA1   4  2 dHDSP_8601
DB1   4 15 dHDSP_8601
DC1   4 13 dHDSP_8601
DD1   4 11 dHDSP_8601
DE1   4  5 dHDSP_8601
DF1   4  3 dHDSP_8601
DG1   4 14 dHDSP_8601
DDP1  4 10 dHDSP_8601

DA2   6  2 dHDSP_8601
DB2   6 15 dHDSP_8601
DC2   6 13 dHDSP_8601
DD2   6 11 dHDSP_8601
DE2   6  5 dHDSP_8601
DF2   6  3 dHDSP_8601
DG2   6 14 dHDSP_8601
DDP2  6 10 dHDSP_8601

DA3  12  2 dHDSP_8601
DB3  12 15 dHDSP_8601
DC3  12 13 dHDSP_8601
DD3  12 11 dHDSP_8601
DE3  12  5 dHDSP_8601
DF3  12  3 dHDSP_8601
DG3  12 14 dHDSP_8601
DDP3 12 10 dHDSP_8601

DA4  17  2 dHDSP_8601
DB4  17 15 dHDSP_8601
DC4  17 13 dHDSP_8601
DD4  17 11 dHDSP_8601
DE4  17  5 dHDSP_8601
DF4  17  3 dHDSP_8601
DG4  17 14 dHDSP_8601
DDP4 17 10 dHDSP_8601

.MODEL dHDSP_8601 D
+ (  
+     IS = 3.97670539E-22 
+      N = 1.67603447 
+     RS = 9.10910000 
+     BV = 50
+    IBV = 100u 
+ )    

.ENDS HDSP_8601
*  
* Diode Model Produced by Altium Ltd  
* Date:  10-Mar-2004 
*  
* Manufacturer: Agilent  
* Component Name: HDSP-513A  
*  
* Parameters derived from information available in data sheet.  
*  
*                 anode-e 
*                 |  anode-d 
*                 |  |  common-cathode 
*                 |  |  |  anode-c 
*                 |  |  |  |  anode-DP 
*                 |  |  |  |  |  anode-b 
*                 |  |  |  |  |  |  anode-a 
*                 |  |  |  |  |  |  |  common-cathode 
*                 |  |  |  |  |  |  |  |  anode-f 
*                 |  |  |  |  |  |  |  |  |  anode-g
*                 |  |  |  |  |  |  |  |  |  |
.SUBCKT HDSP_513A 1  2  3  4  5  6  7  8  9  10

DA1  7 3 dHDSP_513A
DB1  6 3 dHDSP_513A
DC1  4 3 dHDSP_513A
DD1  2 3 dHDSP_513A
DE1  1 3 dHDSP_513A
DF1  9 3 dHDSP_513A
DG1 10 3 dHDSP_513A

DA2  7 8 dHDSP_513A
DB2  6 8 dHDSP_513A
DC2  4 8 dHDSP_513A
DD2  2 8 dHDSP_513A
DE2  1 8 dHDSP_513A
DF2  9 8 dHDSP_513A
DG2 10 8 dHDSP_513A

.MODEL dHDSP_513A D
+ (  
+    IS  = 4.92088043E-22 
+     N  = 1.51994259 
+    RS  = 3.79496255
+    BV  = 4.5
+   IBV  = 100u 
+ )  

.ENDS HDSP_513A
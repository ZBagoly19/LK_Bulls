*  
* Diode Model Produced by Altium Ltd  
* Date:  7-Apr-2004 
*  
* Manufacturer: Agilent  
* Component Name: 5082-7663  
*  
* Parameters derived from information available in data sheet.  
* 
*                 anode-a
*                 |  anode-f
*                 |  |  common-cathode
*                 |  |  |  anode-e
*                 |  |  |  |  anode-d
*                 |  |  |  |  |  anode-DP
*                 |  |  |  |  |  |  anode-c
*                 |  |  |  |  |  |  |  anode-g
*                 |  |  |  |  |  |  |  |  anode-b
*                 |  |  |  |  |  |  |  |  |  common-cathode
*                 |  |  |  |  |  |  |  |  |  |
.SUBCKT 5082_7663 1  2  3  7  8  9  10 11 13 14

DA1   1  3 d5082_7663
DB1  13  3 d5082_7663
DC1  10  3 d5082_7663
DD1   8  3 d5082_7663
DE1   7  3 d5082_7663
DF1   2  3 d5082_7663
DG1  11  3 d5082_7663
DDP1  9  3 d5082_7663

DA2   1 14 d5082_7663
DB2  13 14 d5082_7663
DC2  10 14 d5082_7663
DD2   8 14 d5082_7663
DE2   7 14 d5082_7663
DF2   2 14 d5082_7663
DG2  11 14 d5082_7663
DDP2  9 14 d5082_7663

.MODEL d5082_7663 D
+ (  
+     IS = 6.04055825E-18 
+      N = 1.90788337 
+     RS = 23.52447762 
+     BV = 40
+    IBV = 100u 
+ )  

.ENDS 5082_7663
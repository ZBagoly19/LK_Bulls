*  
* Diode Model Produced by Altium Ltd  
* Date:  10-Mar-2004 
*  
* Manufacturer: Agilent  
* Component Name: HDSP-513E  
*  
* Parameters derived from information available in data sheet.  
*  
*                 anode-e 
*                 |  anode-d 
*                 |  |  common-cathode 
*                 |  |  |  anode-c 
*                 |  |  |  |  anode-DP 
*                 |  |  |  |  |  anode-b 
*                 |  |  |  |  |  |  anode-a 
*                 |  |  |  |  |  |  |  common-cathode 
*                 |  |  |  |  |  |  |  |  anode-f 
*                 |  |  |  |  |  |  |  |  |  anode-g
*                 |  |  |  |  |  |  |  |  |  |
.SUBCKT HDSP_513E 1  2  3  4  5  6  7  8  9  10

DA1  7 3 dHDSP_513E
DB1  6 3 dHDSP_513E
DC1  4 3 dHDSP_513E
DD1  2 3 dHDSP_513E
DE1  1 3 dHDSP_513E
DF1  9 3 dHDSP_513E
DG1 10 3 dHDSP_513E

DA2  7 8 dHDSP_513E
DB2  6 8 dHDSP_513E
DC2  4 8 dHDSP_513E
DD2  2 8 dHDSP_513E
DE2  1 8 dHDSP_513E
DF2  9 8 dHDSP_513E
DG2 10 8 dHDSP_513E

.MODEL dHDSP_513E D
+ (  
+     IS = 6.44208414E-14 
+      N = 2.73863792 
+     RS = 11.58628790 
+     BV = 4.5
+    IBV = 100u 
+ )  

.ENDS HDSP_513E
*  
* Diode Model Produced by Altium Ltd  
* Date:  7-Apr-2004 
*  
* Manufacturer: Agilent  
* Component Name: HDSP-3901  
*  
* Parameters derived from information available in data sheet.  
* 
*                 cathode-a 
*                 |  cathode-f 
*                 |  |  common-anode
*                 |  |  |  cathode-e 
*                 |  |  |  |  common-anode 
*                 |  |  |  |  |  cathode-DP 
*                 |  |  |  |  |  |  cathode-d 
*                 |  |  |  |  |  |  |  common-anode 
*                 |  |  |  |  |  |  |  |  cathode-c 
*                 |  |  |  |  |  |  |  |  |  cathode-g 
*                 |  |  |  |  |  |  |  |  |  |  cathode-b 
*                 |  |  |  |  |  |  |  |  |  |  |  common-anode
*                 |  |  |  |  |  |  |  |  |  |  |  |
.SUBCKT HDSP_3901 2  3  4  5  6  10 11 12 13 14 15 17

DA1   4  2 dHDSP_3901
DB1   4 15 dHDSP_3901
DC1   4 13 dHDSP_3901
DD1   4 11 dHDSP_3901
DE1   4  5 dHDSP_3901
DF1   4  3 dHDSP_3901
DG1   4 14 dHDSP_3901
DDP1  4 10 dHDSP_3901

DA2   6  2 dHDSP_3901
DB2   6 15 dHDSP_3901
DC2   6 13 dHDSP_3901
DD2   6 11 dHDSP_3901
DE2   6  5 dHDSP_3901
DF2   6  3 dHDSP_3901
DG2   6 14 dHDSP_3901
DDP2  6 10 dHDSP_3901

DA3  12  2 dHDSP_3901
DB3  12 15 dHDSP_3901
DC3  12 13 dHDSP_3901
DD3  12 11 dHDSP_3901
DE3  12  5 dHDSP_3901
DF3  12  3 dHDSP_3901
DG3  12 14 dHDSP_3901
DDP3 12 10 dHDSP_3901

DA4  17  2 dHDSP_3901
DB4  17 15 dHDSP_3901
DC4  17 13 dHDSP_3901
DD4  17 11 dHDSP_3901
DE4  17  5 dHDSP_3901
DF4  17  3 dHDSP_3901
DG4  17 14 dHDSP_3901
DDP4 17 10 dHDSP_3901


.MODEL dHDSP_3901 D
+ (  
+     IS = 1E-13 
+      N = 2.7
+     RS = 6.22331865 
+     BV = 2.25
+    IBV = 100u 
+ )  

.ENDS HDSP_3901
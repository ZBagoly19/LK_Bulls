*  
* Diode Model Produced by Altium Ltd  
* Date:  10-Mar-2004 
*  
* Manufacturer: Agilent  
* Component Name: HDSP-H213  
*  
* Parameters derived from information available in data sheet.  
* 
*                 anode-e
*                 |  anode-d
*                 |  |  common-cathode
*                 |  |  |  anode-c
*                 |  |  |  |  anode-DP
*                 |  |  |  |  |  anode-b
*                 |  |  |  |  |  |  anode-a
*                 |  |  |  |  |  |  |  common-cathode
*                 |  |  |  |  |  |  |  |  anode-f
*                 |  |  |  |  |  |  |  |  |  anode-g
*                 |  |  |  |  |  |  |  |  |  | 
.SUBCKT HDSP_H213 1  2  3  4  5  6  7  8  9  10

DA1    7  3  dHDSP_H213
DB1    6  3  dHDSP_H213
DC1    4  3  dHDSP_H213
DD1    2  3  dHDSP_H213
DE1    1  3  dHDSP_H213
DF1    9  3  dHDSP_H213
DG1   10  3  dHDSP_H213
DDP1   5  3  dHDSP_H213

DA2    7  8  dHDSP_H213
DB2    6  8  dHDSP_H213
DC2    4  8  dHDSP_H213
DD2    2  8  dHDSP_H213
DE2    1  8  dHDSP_H213
DF2    9  8  dHDSP_H213
DG2   10  8  dHDSP_H213
DDP2   5  8  dHDSP_H213

.MODEL dHDSP_H213 D
+ (  
+     IS = 2.92097419E-52 
+      N = 0.52799867 
+     RS = 25.27044243 
+     BV = 30
+    IBV = 100u 
+ ) 

.ENDS HDSP_H213